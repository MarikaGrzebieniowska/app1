��;     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.3.0�ub�n_estimators�Kd�estimator_params�(hhhhhhhhhht��base_estimator��
deprecated��	bootstrap���	oob_score���n_jobs�NhK*�verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        hG?�      hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h*�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Pclass��Sex��Age��SibSp��Parch��Fare��Embarked�et�b�n_features_in_�K�
n_outputs_�K�classes_�h)h,K ��h.��R�(KK��h3�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hG?�      hNhJf��_hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h3�f8�����R�(KhLNNNJ����J����K t�b�C              �?�t�bhPh'�scalar���hKC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK�
node_count�Kq�nodes�h)h,K ��h.��R�(KKq��h3�V64�����R�(Kh7N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(h|h3�i8�����R�(KhLNNNJ����J����K t�bK ��h}h�K��h~h�K��hh\K��h�h\K ��h�h�K(��h�h\K0��h�h3�u1�����R�(Kh7NNNJ����J����K t�bK8��uK@KKt�b�B@         P                    �?z����?�           @�@Lq�A�?       E                 �U�R@�x�c���?T           Ȁ@      @       4                    �?��^-��?3           `~@      @                            �?�T�p �?�            @w@       @                          �B@�1�`jg�?"            �K@      @������������������������       ����Q��?             D@       @������������������������       �        	             .@      �?                          �4@��3֞�?�            �s@       @	                        pf� @d}h���?             <@       
                        P�@      �?             0@       ������������������������       ������H�?             "@^      ������������������������       �����X�?             @g      ������������������������       �                     (@>              3                 0C�E@�e!p���?�            r@                                �9@xzY���?�            �q@        ������������������������       �                      G@�                                   @H�f�i��?�            @m@                                   �?`�H�/��?#            �I@        ������������������������       �����X�?             @#                                �7@t��ճC�?             F@                                @D@�7��?            �C@       ������������������������       �                     7@!       ������������������������       �      �?	             0@4       ������������������������       �z�G�z�?             @,                                 �;@(��+�?l            �f@                               pf� @X�<ݚ�?             "@        ������������������������       �      �?             @�       ������������������������       ����Q��?             @�             2                 0#6@�:���?d            �e@             %                   �<@ �Cc}�?`             e@             "                    �?���L��?6            �V@                !                 ���@�����H�?             ;@        ������������������������       �                     $@        ������������������������       �@�0�!��?	             1@        #       $                 �Y5@     �?)             P@        ������������������������       �؇���X�?             5@        ������������������������       �                    �E@        &       +                 �?�@� ���?*            @S@        '       (                    �?@-�_ .�?            �B@        ������������������������       ������H�?             "@        )       *                 �&B@h�����?             <@       ������������������������       �                     3@        ������������������������       ������H�?             "@        ,       /                   @@@      �?             D@        -       .                   �?@      �?             (@        ������������������������       �      �?             @        ������������������������       �      �?             @        0       1                 @3�@؇���X�?             <@        ������������������������       ����Q��?             $@        ������������������������       �        
             2@        ������������������������       ��q�q�?             @        ������������������������       �X�<ݚ�?             "@        5       :                   �;@P����?I            �\@        6       9                   �7@�p����?#            �N@       7       8                    �?��B����?             J@       ������������������������       �*O���?             B@        ������������������������       �      �?             0@        ������������������������       �                     "@        ;       >                     @�T`�[k�?&            �J@        <       =                   �H@`2U0*��?             9@     �?������������������������       �                     5@      �?������������������������       �      �?             @      �??       @                 �̌@��>4և�?             <@      �?������������������������       �"pc�
�?             &@      �?A       B                    �?��.k���?             1@      �?������������������������       �      �?             @      �?C       D                 @3#%@��
ц��?
             *@      �?������������������������       �                     @      �?������������������������       �      �?              @      �?F       K                   �A@>a�����?!            �I@     �?G       J                    �?l��\��?             A@     �?H       I                 �_@��2(&�?
             6@      �?������������������������       ���S�ۿ?             .@      �?������������������������       �����X�?             @      �?������������������������       �        	             (@      �?L       O                   �G@�t����?             1@     �?M       N                   @D@���Q��?             $@      �?������������������������       ��q�q�?             @      �?������������������������       �      �?             @      �?������������������������       �؇���X�?             @      �?Q       R                    �?s8?U��?o            �e@      �?������������������������       ������H�?             "@      �?S       ^                    �?��a����?i            �d@      �?T       U                    0@��G���?0            �R@      �?������������������������       �      �?             (@      �?V       W                    @��� ��?)             O@      �?������������������������       �և���X�?             @      �?X       Y                    �?,�+�C�?$            �K@      �?������������������������       �      �?              @      �?Z       [                   `B@`Ql�R�?            �G@     �?������������������������       �                     A@      �?\       ]                    H@$�q-�?	             *@      �?������������������������       �؇���X�?             @      �?������������������������       �                     @        _       f                    �?�5��
J�?9             W@        `       e                 м�9@��0{9�?            �G@        a       d                   �>@�X����?             6@       b       c                    �?��S���?
             .@        ������������������������       �      �?              @        ������������������������       �����X�?             @        ������������������������       �                     @        ������������������������       �                     9@        g       h                    �?�q�q�?            �F@        ������������������������       �                     @        i       p                   �=@�n_Y�K�?            �C@       j       k                    �?X�<ݚ�?             ;@        ������������������������       �                     @       l       o                    @�X����?             6@       m       n                     @���Q��?	             .@       ������������������������       �      �?              @       ������������������������       �                     @        ������������������������       �؇���X�?             @        ������������������������       �                     (@       �t�b�values�h)h,K ��h.��R�(KKqKK��h\�B       �{@     �p@     �v@     �e@     @v@     @`@     �s@     �K@     �C@      0@      8@      0@      .@             `q@     �C@      6@      @      $@      @       @      �?       @      @      (@              p@     �@@     `o@      =@      G@             �i@      =@      G@      @      @       @     �D@      @     �B@       @      7@              ,@       @      @      �?     �c@      8@      @      @       @       @      @       @     @c@      4@     �b@      2@     @U@      @      8@      @      $@              ,@      @     �N@      @      2@      @     �E@             @P@      (@     �A@       @       @      �?      ;@      �?      3@               @      �?      >@      $@      @      @      @      @      @      @      8@      @      @      @      2@              @       @      @      @     �C@     �R@      ;@      A@      ;@      9@      *@      7@      ,@       @              "@      (@     �D@      �?      8@              5@      �?      @      &@      1@       @      "@      "@       @       @       @      @      @      @               @      @       @     �E@      @      ?@      @      3@      �?      ,@       @      @              (@      @      (@      @      @       @      @       @       @      �?      @     �T@      W@      �?       @     �T@      U@      N@      ,@      @      @      K@       @      @      @     �I@      @      @      @      G@      �?      A@              (@      �?      @      �?      @              6@     �Q@      @      D@      @      .@      @       @       @      @      @       @              @              9@      .@      >@              @      .@      8@      .@      (@              @      .@      @      "@      @       @      @      @              @      �?              (@�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�=�KhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK	hsKKhth)h,K ��h.��R�(KKK��h{�B�         &                    �?��!h
��?�           @�@Lq�A�?                            �?tk~X��?           @}@ �=	�                            �G@#z�i��?0            �T@�@	�                           x#J@�&�5y�?$             O@ �h��                             =@��hJ,�?             A@ ,]qG�?������������������������       �����X�?             ,@��yr�J�������������������������       �P���Q�?             4@�&g��v0                           �?և���X�?             <@ �����	       
                   �;@���Q��?	             .@ܹ:�B5������������������������       �      �?              @~����,�������������������������       �����X�?             @a                              03U@��
ц��?
             *@        ������������������������       �����X�?             @�       ������������������������       ��q�q�?             @f                                  @@�G�z��?             4@        ������������������������       �z�G�z�?             @                                 �K@��S���?             .@        ������������������������       �      �?              @       ������������������������       �և���X�?             @#                                 $@$�D�B{�?�             x@                                  @�q�q�?             5@       ������������������������       �                     *@!       ������������������������       �      �?              @4              %                    �?H��g���?�            �v@              $                 0�_F@V1��=��?�            �r@                                 �?��o�um�?�            0r@        ������������������������       ��t����?             A@�              !                    �?edc�?�            p@                                ��@�����H�?             B@       ������������������������       �                     "@�                                 �=@PN��T'�?             ;@       ������������������������       �z�G�z�?
             4@�       ������������������������       �                     @�      "       #                 ��@�;��?�            �k@        ������������������������       ���Y��]�?            �D@�      ������������������������       �DG��L�?t            �f@�       ������������������������       �r�q��?             @[      ������������������������       �        %             Q@/      '       4                     @�Ee@���?�            �n@      (       1                  "�b@      �?Y             `@      )       0                   �H@����q�?O            @[@      *       /                   �;@�a�O�?F            @X@       +       .                    �?��Y��]�?            �D@        ,       -                   �7@�}�+r��?             3@       ������������������������       �z�G�z�?             @        ������������������������       �        
             ,@        ������������������������       �                     6@        ������������������������       �        )             L@        ������������������������       ��8��8��?	             (@        2       3                    :@�KM�]�?
             3@        ������������������������       �����X�?             @        ������������������������       �                     (@        5       H                 03�7@�'�ſ:�?L             ]@       6       C                 ��.@0d4�[%�?>            �W@       7       >                   �9@���Q��?+            @P@        8       =                    �?��S���?             >@       9       :                    �?���Q��?             9@        ������������������������       ��q�q�?             @        ;       <                   �5@D�n�3�?             3@        ������������������������       �      �?              @        ������������������������       ����|���?             &@        ������������������������       �z�G�z�?             @        ?       B                    �?����X�?            �A@       @       A                    �?�n`���?             ?@       ������������������������       ��<ݚ�?             2@        ������������������������       �8�Z$���?             *@        ������������������������       �                     @        D       E                    �?ףp=
�?             >@        ������������������������       �                     *@        F       G                 pff0@@�0�!��?             1@        ������������������������       ��<ݚ�?             "@        ������������������������       �      �?              @        I       J                 ��T?@���N8�?             5@       ������������������������       �        	             .@        ������������������������       �r�q��?             @        �t�bh�h)h,K ��h.��R�(KKKKK��h\�B�       �z@     �q@     �w@     �V@      K@      <@     �F@      1@      =@      @      $@      @      3@      �?      0@      (@      "@      @      @      @      @       @      @      @      @       @       @      @      "@      &@      �?      @       @      @      @      @      @      @     0t@     �O@      @      ,@              *@      @      �?     �s@     �H@      o@     �H@     �n@      F@      8@      $@     �k@      A@      @@      @      "@              7@      @      0@      @      @             �g@      >@      D@      �?     �b@      =@      �?      @      Q@             �J@     �g@      @      _@       @     �Z@      �?      X@      �?      D@      �?      2@      �?      @              ,@              6@              L@      �?      &@       @      1@       @      @              (@     �H@     �P@      =@     �P@      :@     �C@      0@      ,@      .@      $@      @       @      &@       @      @      @      @      @      �?      @      $@      9@      @      9@      @      ,@       @      &@      @              @      ;@              *@      @      ,@       @      @      �?      @      4@      �?      .@              @      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ\bshG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK
hsKghth)h,K ��h.��R�(KKg��h{�B�         0                     @z��Y�)�?�           @�@ Lq�A�?                          �,@�G��l��?�            �s@      (@                           �?PN���?8            @V@ �B	�  ������������������������       �                      @��?	�                             �?ڤ���?3            @T@    �O@                           @     p�?(             P@     �H@������������������������       �                     &@      A@                          �F@0��_��?!            �J@     @	                          �;@X�EQ]N�?            �E@     =@
                           &@�>����?             ;@      _@������������������������       �      �?              @      2@������������������������       �        
             3@      L@                          �'@     ��?             0@        ������������������������       �                     @      ,@������������������������       ��q�q�?             "@      @������������������������       �                     $@      9@������������������������       ��t����?             1@               /                   �M@��^w��?�            @l@              "                    �?4C)�m��?�            @k@                                   &@�*/�8V�?@            �W@        ������������������������       �                     &@                                   �?�1/z��?9            �T@                               ��$:@     ��?-             P@        ������������������������       �                     $@                                   �?�<ݚ�?&             K@      �?������������������������       �      �?             0@      �?                          �G@���y4F�?             C@     �?                            �?�>����?             ;@     �?������������������������       ��C��2(�?             6@      �?������������������������       �                     @      �?������������������������       ��eP*L��?             &@      �?        !                    �?�}�+r��?             3@      �?������������������������       �      �?              @3      ������������������������       �                     &@A      #       ,                  "�b@�7���?E             _@       $       '                   �;@` A�c̭?9             Y@        %       &                    :@`Jj��?             ?@        ������������������������       �      �?              @j       ������������������������       �                     7@�       (       +                    �?@	tbA@�?&            @Q@        )       *                 �U5Q@�IєX�?
             1@        ������������������������       �؇���X�?             @�       ������������������������       �                     $@$       ������������������������       �                     J@       -       .                 `D�c@�q�q�?             8@        ������������������������       �և���X�?             ,@-       ������������������������       �                     $@]       ������������������������       �                      @�       1       R                    �?7����?�            �x@       2       A                 �?�@����?�            pq@        3       @                 �1@X�GP>��?V            �_@       4       ?                 ��@����\�?>            �V@       5       :                   �:@ �\���?7            �S@        6       9                    7@      �?             8@      7       8                 �Y�@      �?             0@        ������������������������       �                     "@`      ������������������������       �؇���X�?             @:      ������������������������       �      �?              @;      ;       >                    �? �Jj�G�?$            �K@       <       =                 ���@��S�ۿ?             .@      ������������������������       �                     $@7      ������������������������       �z�G�z�?             @G       ������������������������       �                     D@      ������������������������       ����!pc�?             &@!      ������������������������       �                    �B@�      B       C                    �?$�Z����?\             c@       ������������������������       �      �?             (@8       D       I                    $@(N:!���?V            �a@       E       H                    @      �?             4@      F       G                    @�z�G��?             $@       ������������������������       �z�G�z�?             @,      ������������������������       ����Q��?             @�      ������������������������       �z�G�z�?             $@�       J       K                 @3�@�.�?�P�?H             ^@        ������������������������       �����X�?             @v      L       O                    �?ЮN
��?B            @\@      M       N                 ���#@ �q�q�?8             X@      ������������������������       � 	��p�?$             M@�      ������������������������       �                     C@�      P       Q                    ;@�t����?
             1@       ������������������������       �                     @�       ������������������������       �r�q��?             (@      S       b                 03�7@�ݜ����?G            �]@      T       U                    @      �?6             V@       ������������������������       ������H�?             "@g      V       W                   �5@�����?1            �S@        ������������������������       ��ՙ/�?             5@y       X       Y                 �̌@T����1�?$             M@        ������������������������       �                     0@�       Z       [                    �?��6���?             E@        ������������������������       ������H�?             "@        \       ]                 @3�@�eP*L��?            �@@        ������������������������       �����X�?             @        ^       a                   �=@�n_Y�K�?             :@       _       `                   �.@      �?	             (@        ������������������������       �                     @        ������������������������       �և���X�?             @        ������������������������       �      �?             ,@        c       f                 ��p@@(;L]n�?             >@       d       e                    @@4և���?
             ,@        ������������������������       �z�G�z�?             @        ������������������������       �                     "@        ������������������������       �                     0@        �t�bh�h)h,K ��h.��R�(KKgKK��h\�Bp       �|@     @o@     �b@     �d@     �N@      <@               @     �N@      4@     �M@      @      &@              H@      @      C@      @      9@       @      @       @      3@              *@      @      @              @      @      $@               @      .@     @V@      a@     @T@      a@     �Q@      8@              &@     �Q@      *@      J@      (@      $@              E@      (@      (@      @      >@       @      9@       @      4@       @      @              @      @      2@      �?      @      �?      &@              &@     @\@      @     @X@       @      =@       @      @              7@      �?      Q@      �?      0@      �?      @              $@              J@       @      0@       @      @              $@       @             �s@     @U@     @o@      =@      ^@      @     �T@      @     �R@      @      5@      @      .@      �?      "@              @      �?      @       @      K@      �?      ,@      �?      $@              @      �?      D@               @      @     �B@             @`@      6@      @      @      _@      0@      .@      @      @      @      @      �?      @       @       @       @     @[@      &@       @      @     �Z@      @      W@      @      K@      @      C@              .@       @      @              $@       @      O@      L@     �@@     �K@      �?       @      @@     �G@      *@       @      3@     �C@              0@      3@      7@      �?       @      2@      .@       @      @      0@      $@      "@      @      @              @      @      @      @      =@      �?      *@      �?      @      �?      "@              0@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��.hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKmhth)h,K ��h.��R�(KKm��h{�B@         J                    �?��!h
��?�           @�@      @                           @�՘���?'           �}@                                   @�q�q�?            �@@0��  ������������������������       �                     4@�����  ������������������������       �8�Z$���?             *@      8@                          �8@�t�i�?           �{@                                   �?�ڊ�e��?=             Y@      @                            @ ,U,?��?3            �T@      �?	       
                    4@���7�?             6@    @X@������������������������       �ףp=
�?             $@      Q@������������������������       �                     (@      J@                           �?��GEI_�?&            �N@        ������������������������       �և���X�?             @�                               @3�@@3����?!             K@        ������������������������       �                     9@      �?                          �3@XB���?             =@      @������������������������       ������H�?             "@        ������������������������       �                     4@  �@  �?                           �?������?
             1@ ��@���@������������������������       �      �?             @        ������������������������       ��C��2(�?             &@               9                 ���=@�YC�ż�?�            `u@̀A�̀A       ,                   @@@Rq�����?�            �o@ �A  �A                           �?     ��?e             d@                                ���@f���M�?             ?@        ������������������������       �                     @gD(AfffA������������������������       �� �	��?             9@  �?  �?                            @&^�)b�?R             `@       @������������������������       ��8��8��?             8@       @                           �?�϶O'3�?E            @Z@       @������������������������       ��㙢�c�?             7@       @        #                   �;@��P���?7            �T@       @!       "                 ��L@X�<ݚ�?             2@      ������������������������       ����|���?             &@A      ������������������������       �؇���X�?             @�       $       +                   �>@     ��?*             P@       %       *                    �?h�WH��?$             K@       &       )                 ��) @�����H�?            �F@       '       (                 �?$@�g�y��?             ?@        ������������������������       �؇���X�?             @�       ������������������������       �                     8@�       ������������������������       �����X�?             ,@�       ������������������������       �                     "@$       ������������������������       �      �?             $@       -       0                     �?<����?<            �W@        .       /                   �G@���y4F�?             3@       ������������������������       �$�q-�?             *@]       ������������������������       �      �?             @�       1       6                   �E@�}�+r��?1             S@       2       5                    �? pƵHP�?             J@       3       4                 `fF)@P�Lt�<�?             C@       ������������������������       �                     ?@�       ������������������������       �؇���X�?             @�       ������������������������       �                     ,@      7       8                   �'@      �?             8@       ������������������������       �z�G�z�?             .@`      ������������������������       �                     "@:      :       ;                   �>@�f7�z�?6            �U@       ������������������������       �8�Z$���?             *@?      <       ?                  x#J@~�hP��?.            �R@       =       >                   �B@���7�?             6@       ������������������������       �؇���X�?             @G       ������������������������       �        	             .@      @       C                    �?��
ц��?              J@       A       B                 ��+T@�����?             3@       ������������������������       ��<ݚ�?             "@�      ������������������������       ����Q��?             $@8       D       I                    �?�q�q�?            �@@      E       F                 `�jM@
j*D>�?             :@       ������������������������       �����X�?             ,@-      G       H                   �H@�8��8��?             (@       ������������������������       �z�G�z�?             @�      ������������������������       �                     @�       ������������������������       �                     @�       K       T                 `f�$@N��6z�?�            �m@       L       O                   �9@�g�y��?"             O@       M       N                   �1@X�Cc�?             <@       ������������������������       ��q�q�?             "@�      ������������������������       ����y4F�?             3@�      P       Q                    �?j���� �?             A@       ������������������������       ������?	             3@�       R       S                    >@��S���?	             .@      ������������������������       ��q�q�?             "@-      ������������������������       ��q�q�?             @%      U       d                     @ �ܽ��?r            �e@      V       a                   �H@H�Swe�?R            @_@       W       ^                 ���a@Ц�f*�?G            �[@       X       ]                    6@�L��ȕ?<            @W@        Y       Z                    �?(;L]n�?             >@        ������������������������       �                     "@        [       \                    ?@���N8�?             5@        ������������������������       ������H�?             "@        ������������������������       �                     (@        ������������������������       �        +            �O@        _       `                    �?�t����?             1@       ������������������������       �                     (@        ������������������������       ����Q��?             @        b       c                   �I@z�G�z�?             .@        ������������������������       �      �?             @        ������������������������       �                     "@        e       j                 ���4@z�):���?              I@        f       i                   �=@������?             >@       g       h                    �?�㙢�c�?             7@        ������������������������       ��	j*D�?             *@        ������������������������       �                     $@        ������������������������       �և���X�?             @        k       l                    #@P���Q�?             4@        ������������������������       �      �?             @        ������������������������       �                     0@        �t�bh�h)h,K ��h.��R�(KKmKK��h\�B�       �z@     �q@     �v@     �[@      &@      6@              4@      &@       @      v@      V@     �V@      "@     �S@      @      5@      �?      "@      �?      (@             �L@      @      @      @     �J@      �?      9@              <@      �?       @      �?      4@              *@      @      @      @      $@      �?     pp@     �S@     �j@     �E@     @_@     �A@      4@      &@      @              ,@      &@     @Z@      8@      6@       @     �T@      6@      3@      @      P@      2@      $@       @      @      @      @      �?      K@      $@     �H@      @      D@      @      >@      �?      @      �?      8@              $@      @      "@              @      @     �U@       @      .@      @      (@      �?      @      @      R@      @     �I@      �?     �B@      �?      ?@              @      �?      ,@              5@      @      (@      @      "@             �I@      B@       @      &@     �H@      9@      5@      �?      @      �?      .@              <@      8@      @      *@       @      @      @      @      6@      &@      .@      &@      @      $@      &@      �?      @      �?      @              @             @P@     �e@      @@      >@      2@      $@      @      @      .@      @      ,@      4@      @      *@       @      @      @      @       @      @     �@@     �a@      @     �]@      @     �Z@      �?      W@      �?      =@              "@      �?      4@      �?       @              (@             �O@       @      .@              (@       @      @      @      (@      @      @              "@      ;@      7@       @      6@      @      3@      @      "@              $@      @      @      3@      �?      @      �?      0@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJj�c;hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKwhth)h,K ��h.��R�(KKw��h{�B�         L                    �?�)�>_M�?�           @�@      @                           $@�g[Z��?            P|@ TC��                            �;@և���X�?             <@ A	�  ������������������������       �                     $@�) 	�                             @�q�q�?             2@      @������������������������       �                     @     �A@������������������������       �$�q-�?             *@      8@                           �?���f_�?           �z@      2@	                            �?�	j*D�?2            �S@      $@
                        ��hU@���>4��?             <@     �?                           A@�eP*L��?             6@     @                        ��>@�n_Y�K�?	             *@      @������������������������       �      �?             @�       ������������������������       �����X�?             @      @������������������������       ��<ݚ�?             "@      9@������������������������       �r�q��?             @      8@                        83##@j�q����?              I@                              ���@�C��2(�?            �@@       ������������������������       �                     *@�      ������������������������       �R���Q�?             4@w                                  @ҳ�wY;�?             1@       ������������������������       �      �?              @�      ������������������������       �X�<ݚ�?             "@�             7                   �<@�-q���?�            �u@             2                 `fF:@���(ͷ�?�            `i@             +                    �?����?o            �e@                                 �?�X�<ݺ?\             b@                                ��@      �?             0@       ������������������������       �                     @�      ������������������������       ��C��2(�?             &@(                                  1@     x�?Q             `@       ������������������������       �      �?              @J      !       (                 �1@(;L]n�?K             ^@       "       #                 `f�@l��\��?             A@       ������������������������       �                     &@�       $       %                 ���@�LQ�1	�?             7@        ������������������������       ��q�q�?             @v       &       '                    7@�IєX�?             1@        ������������������������       �r�q��?             @�       ������������������������       �                     &@�       )       *                   �;@��f�{��?5            �U@       ������������������������       �                    �F@�       ������������������������       ���Y��]�?            �D@$       ,       1                    �?z�G�z�?             >@       -       0                   �9@��<b���?             7@       .       /                    5@�n_Y�K�?             *@        ������������������������       ��q�q�?             @]       ������������������������       �և���X�?             @�       ������������������������       �                     $@A       ������������������������       �؇���X�?             @�       3       4                   �>@д>��C�?             =@        ������������������������       �      �?             @�       5       6                    �?HP�s��?             9@       ������������������������       �؇���X�?             ,@      ������������������������       �                     &@�       8       C                   @E@8��8���?X             b@      9       B                   �D@�4���L�?3            �U@      :       A                 0�K@� ���?.            @S@      ;       >                   @@@���Ls�?)            @P@       <       =                     @д>��C�?             =@       ������������������������       �                     @7      ������������������������       ���<b���?             7@G       ?       @                 03�3@������?             B@      ������������������������       �                     =@!      ������������������������       �؇���X�?             @�      ������������������������       �      �?             (@�      ������������������������       �X�<ݚ�?             "@8       D       G                 `fF:@ 	��p�?%             M@      E       F                   @L@��Y��]�?            �D@      ������������������������       �                     A@-      ������������������������       �؇���X�?             @,      H       K                    L@@�0�!��?             1@      I       J                 �T!@@�z�G��?
             $@        ������������������������       �      �?             @�       ������������������������       �                     @v      ������������������������       �                     @�      M       \                     @�T����?�            0p@      N       Y                  "�b@��*����?V            `a@      O       X                    �? _�@�Y�?K             ]@      P       S                    �? ���J��?5            �S@       Q       R                   �H@ 7���B�?             ;@       ������������������������       �                     3@      ������������������������       �      �?              @-      T       W                  �v7@���J��?"            �I@       U       V                    =@�nkK�?             7@       ������������������������       ��C��2(�?             &@�       ������������������������       �        	             (@y       ������������������������       �                     <@}       ������������������������       �                     C@�       Z       [                    �?���}<S�?             7@       ������������������������       �                     0@        ������������������������       �����X�?             @        ]       v                 ��Y7@��0u���?L             ^@       ^       u                   @B@ڡR����?=            �X@       _       d                 ��@�L�lRT�?9            �V@        `       c                    �?�C��2(�?             6@       a       b                  s�@؇���X�?	             ,@       ������������������������       �      �?              @        ������������������������       �r�q��?             @        ������������������������       �                      @        e       j                 `f�%@�ʻ����?,             Q@        f       g                    �?�LQ�1	�?             7@        ������������������������       �؇���X�?             @        h       i                 @33"@      �?             0@       ������������������������       �                     $@        ������������������������       ��q�q�?             @        k       n                    5@�q�q�?            �F@        l       m                    @��.k���?             1@       ������������������������       ������H�?             "@        ������������������������       �                      @        o       t                    �?d}h���?             <@       p       q                    �?�����?             5@        ������������������������       �                      @        r       s                   �>@8�Z$���?             *@        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �և���X�?             @        ������������������������       �                      @        ������������������������       ����7�?             6@        �t�bh�h)h,K ��h.��R�(KKwKK��h\�Bp       `{@      q@     Pw@      T@      (@      0@              $@      (@      @              @      (@      �?     �v@      P@      K@      8@      *@      .@      (@      $@      @       @      @      @       @      @      @       @      �?      @     �D@      "@      >@      @      *@              1@      @      &@      @      @      �?      @      @     0s@      D@      g@      3@      d@      ,@      a@       @      .@      �?      @              $@      �?     @^@      @      @      @      ]@      @      ?@      @      &@              4@      @      @       @      0@      �?      @      �?      &@             @U@      �?     �F@              D@      �?      8@      @      2@      @       @      @      @       @      @      @      $@              @      �?      8@      @      �?      @      7@       @      (@       @      &@             �^@      5@     @Q@      1@     @P@      (@     �M@      @      8@      @      @              2@      @     �A@      �?      =@              @      �?      @      @      @      @      K@      @      D@      �?      A@              @      �?      ,@      @      @      @      �?      @      @              @             @P@     @h@      @     �`@       @     �\@       @      S@      �?      :@              3@      �?      @      �?      I@      �?      6@      �?      $@              (@              <@              C@       @      5@              0@       @      @     �N@     �M@      D@      M@      @@      M@       @      4@       @      (@      �?      @      �?      @               @      >@      C@      .@       @      �?      @      ,@       @      $@              @       @      .@      >@      "@       @      �?       @       @              @      6@       @      3@               @       @      &@              @       @      @      @      @       @              5@      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJGԙGhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKkhth)h,K ��h.��R�(KKk��h{�B�         6                     @�3�n��?�           @�@       @       )                    �?z�J��?�            �t@     P@                           $@J������?�            �h@       @������������������������       �                     @      @                           �??���?{            �g@      @                           �?\�Uo��?             C@     D@       
                    ?@���>4��?             <@     �?       	                   �;@p�ݯ��?             3@      @������������������������       �      �?             @      @������������������������       ��	j*D�?             *@        ������������������������       ��q�q�?             "@      @������������������������       �z�G�z�?             $@      @       (                    �?L紂P�?a             c@                                   �?tK���:�?T            ``@      5@                           �?      �?$             J@     @                           @@      �?             F@                                 �D@��}*_��?             ;@                              ��$:@������?             .@      ������������������������       �                     "@�      ������������������������       ��q�q�?             @w                                �I@      �?	             (@      ������������������������       �և���X�?             @�      ������������������������       ����Q��?             @�                                �=@�IєX�?
             1@      ������������������������       ������H�?             "@�      ������������������������       �                      @c      ������������������������       �      �?              @             #                   �*@$��$�L�?0            �S@                               `f�)@8��8���?             H@                                �E@      �?             @@      ������������������������       � 7���B�?             ;@V      ������������������������       �z�G�z�?             @J      !       "                   �:@     ��?             0@       ������������������������       �                     @A      ������������������������       ��eP*L��?             &@�       $       '                   �@@�g�y��?             ?@        %       &                    �?�8��8��?	             (@        ������������������������       �                     @j       ������������������������       �؇���X�?             @�       ������������������������       �        
             3@�       ������������������������       �                     6@�       *       1                   �;@DgV`�?Q            ``@        +       .                   �7@�C��2(�?#            �K@       ,       -                 83�`@г�wY;�?             A@       ������������������������       �                     >@       ������������������������       �      �?             @-       /       0                    �?��s����?             5@        ������������������������       ����!pc�?             &@�       ������������������������       �ףp=
�?             $@A       2       5                     �?�"w����?.             S@       3       4                   �J@��Y��]�?            �D@        ������������������������       �z�G�z�?             @�       ������������������������       �                     B@�       ������������������������       �                    �A@      7       B                    �?�E�_�?�            �w@        8       =                    �?�qs�_�?E            �Z@      9       :                    �?Z���c��?(            �O@      ������������������������       �p9W��S�?             C@;      ;       <                    �?HP�s��?             9@      ������������������������       �                     1@I      ������������������������       �      �?              @7      >       A                 ��.@      �?             F@       ?       @                    �?�!���?             A@      ������������������������       �����X�?             <@!      ������������������������       �      �?             @�      ������������������������       �                     $@�      C       D                 �ٝ@��X���?�            @q@        ������������������������       �                     @@8      E       X                    �?��f/w�?�            �n@      F       W                    �?ghډC�?c            �b@      G       H                   �0@p^H�&m�?W            �`@       ������������������������       ��q�q�?             @�      I       V                 �T�E@     �?R             `@       J       Q                    ?@��a��?N            @^@       K       L                 �&B@�zvܰ?4             V@       ������������������������       �      �?              @�      M       N                 pf� @@�z�G�?/             T@      ������������������������       �                    �F@�      O       P                 ���!@��?^�k�?            �A@       ������������������������       ������H�?             "@�      ������������������������       �                     :@�       R       S                   @@@<���D�?            �@@       ������������������������       �      �?              @-      T       U                   �E@`2U0*��?             9@      ������������������������       �                     0@g      ������������������������       ������H�?             "@�       ������������������������       �և���X�?             @y       ������������������������       �                     0@}       Y       d                    �?�ހ��?9            �W@       Z       [                 �&B@~|z����?            �J@        ������������������������       �r�q��?             @        \       c                 ��&@z�J��?            �G@       ]       `                   �9@��J�fj�?            �B@        ^       _                   �5@      �?             0@        ������������������������       ��<ݚ�?             "@        ������������������������       �                     @        a       b                   �=@�q�q�?	             5@       ������������������������       ��	j*D�?             *@        ������������������������       �      �?              @        ������������������������       ��z�G��?             $@        e       h                 ���4@���� �?            �D@        f       g                   �*@r�q��?
             (@       ������������������������       �      �?              @        ������������������������       �      �?             @        i       j                    @XB���?             =@        ������������������������       �z�G�z�?             @        ������������������������       �                     8@        �t�bh�h)h,K ��h.��R�(KKkKK��h\�B�       �{@     �p@      d@      e@     `c@     �E@              @     `c@      B@      7@      .@      .@      *@      (@      @      @      @      "@      @      @      @       @       @     �`@      5@     �[@      5@     �C@      *@     �@@      &@      1@      $@      &@      @      "@               @      @      @      @      @      @      @       @      0@      �?       @      �?       @              @       @     �Q@       @     �D@      @      >@       @      :@      �?      @      �?      &@      @      @              @      @      >@      �?      &@      �?      @              @      �?      3@              6@              @     @_@      @      I@      �?     �@@              >@      �?      @      @      1@      @       @      �?      "@      �?     �R@      �?      D@      �?      @              B@             �A@     �q@     �X@     �N@      G@      I@      *@      ;@      &@      7@       @      1@              @       @      &@     �@@      &@      7@       @      4@      @      @              $@      l@      J@      @@              h@      J@      a@      *@     @^@      *@      @       @     @]@      &@     �\@      @     @U@      @      @       @     �S@      �?     �F@              A@      �?       @      �?      :@              =@      @      @      @      8@      �?      0@               @      �?      @      @      0@             �K@     �C@      9@      <@      �?      @      8@      7@      5@      0@      ,@       @      @       @      @              @      ,@      @      "@      @      @      @      @      >@      &@       @      $@      �?      @      �?      @      <@      �?      @      �?      8@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��AhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKqhth)h,K ��h.��R�(KKq��h{�B@         N                    �?ƈ�VM�?�           @�@      @                            �?�����?           �{@      @                          �;@�x_F-�?;            �Y@       @                          �8@     ��?	             0@     &@������������������������       ��<ݚ�?             "@      @������������������������       �                     @      �?                           �?�%^�?2            �U@      @                          �>@      �?"             N@     �?	       
                    �?����"�?             =@      �?������������������������       �      �?             @                                ��$:@���Q��?             9@     �@@������������������������       �                     @       @                          �I@X�<ݚ�?
             2@       ������������������������       �z�G�z�?             $@      G@������������������������       �      �?              @                                `�I@��� ��?             ?@     4@                          �A@���N8�?             5@       ������������������������       �                     (@�      ������������������������       ������H�?             "@�      ������������������������       ��z�G��?             $@w                                 �?R�}e�.�?             :@       ������������������������       �X�<ݚ�?             "@�      ������������������������       �@�0�!��?             1@�                                 @h!�'nf�?�            0u@                                   @�S����?             3@      ������������������������       �                     &@c      ������������������������       �      �?              @             %                     @أp=
��?�             t@              $                    �?�ӖF2��?+            �Q@             #                   @A@l�b�G��?$            �L@                                 �(@������?            �B@       ������������������������       �        	             ,@J      !       "                    �?�㙢�c�?             7@      ������������������������       �@�0�!��?
             1@A      ������������������������       �r�q��?             @�       ������������������������       �                     4@�       ������������������������       �@4և���?             ,@v       &       M                 �T�I@� ��?�             o@       '       *                 ��@\���(\�?�             n@        (       )                 ���@     ��?
             0@        ������������������������       �����X�?             @�       ������������������������       ��q�q�?             "@�       +       J                    0@      �?�             l@       ,       I                    �?(4w%��?y            �g@       -       2                    �?��աU�?s            �f@        .       1                  ��@��G���?            �B@       /       0                 ���@ףp=
�?             4@        ������������������������       ������H�?             "@�       ������������������������       ��C��2(�?             &@A       ������������������������       ��t����?
             1@�       3       <                 �?�@��1���?\             b@       4       7                   �8@(�5�f��?/            �S@        5       6                   �4@�KM�]�?             3@        ������������������������       �                     @      ������������������������       �r�q��?             (@�       8       9                 ��L@ �.�?Ƞ?#             N@       ������������������������       �                     ?@:      :       ;                    ?@XB���?             =@      ������������������������       �                     5@?      ������������������������       �      �?              @I      =       H                   �@@�GN�z�?-            �P@      >       E                 ���!@�E��ӭ�?&             K@       ?       @                   �3@     ��?             @@       ������������������������       ��q�q�?             @!      A       B                   �:@R�}e�.�?             :@       ������������������������       �                      @�      C       D                   �>@b�2�tk�?             2@       ������������������������       ��	j*D�?	             *@8      ������������������������       ����Q��?             @      F       G                    :@"pc�
�?             6@      ������������������������       ��C��2(�?             &@,      ������������������������       ����!pc�?             &@�      ������������������������       �                     (@�       ������������������������       ��<ݚ�?             "@�       K       L                    �?Pa�	�?            �@@       ������������������������       ��C��2(�?             &@�      ������������������������       �                     6@�      ������������������������       �X�<ݚ�?             "@�      O       X                     @2�K^V�?�            �p@      P       U                 ���a@��?^�k�?\            �a@      Q       T                    �? _�@�Y�?O             ]@        R       S                   @H@�FVQ&�?            �@@      ������������������������       �                     <@-      ������������������������       ����Q��?             @%      ������������������������       �        7            �T@g      V       W                 `D�g@�8��8��?             8@        ������������������������       �����X�?             @y       ������������������������       �                     1@}       Y       ^                    �?���nU��?M            ``@        Z       ]                   �8@>��C��?            �E@        [       \                 P��+@��Q��?
             4@       ������������������������       �"pc�
�?             &@        ������������������������       �X�<ݚ�?             "@        ������������������������       ��LQ�1	�?             7@        _       p                    B@7�A�0�?5             V@       `       o                    =@�;�vv��?.            @R@       a       b                 �&B@B�
k���?*            �P@        ������������������������       �r�q��?             (@        c       l                 �̼6@���Q��?$            �K@       d       i                    �?�G��l��?             E@       e       h                 �]*@�q�q�?             >@       f       g                 @3�@���y4F�?             3@        ������������������������       �X�<ݚ�?             "@        ������������������������       �                     $@        ������������������������       ��eP*L��?             &@        j       k                 ���'@r�q��?             (@        ������������������������       �؇���X�?             @        ������������������������       �z�G�z�?             @        m       n                    @8�Z$���?	             *@        ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �r�q��?             @        ������������������������       �                     .@        �t�bh�h)h,K ��h.��R�(KKqKK��h\�B        z@     �r@     �u@     �V@     �Q@      ?@      @      "@      @       @              @      P@      6@     �F@      .@      2@      &@      @      �?      .@      $@      @               @      $@       @       @      @       @      ;@      @      4@      �?      (@               @      �?      @      @      3@      @      @      @      ,@      @     �q@     �M@      @      0@              &@      @      @     Pq@     �E@     �P@      @     �J@      @     �@@      @      ,@              3@      @      ,@      @      @      �?      4@              *@      �?     `j@      C@     �i@     �@@      &@      @      @       @      @      @     �h@      <@     �d@      ;@     �c@      9@      >@      @      2@       @       @      �?      $@      �?      (@      @     �_@      2@      S@      @      1@       @      @              $@       @     �M@      �?      ?@              <@      �?      5@              @      �?     �I@      .@     �C@      .@      5@      &@       @      @      3@      @       @              &@      @      "@      @       @      @      2@      @      $@      �?       @      @      (@              @       @      @@      �?      $@      �?      6@              @      @     @P@     �i@      @      a@       @     �\@       @      ?@              <@       @      @             �T@       @      6@       @      @              1@     �N@     �Q@      $@     �@@      @      *@       @      "@      @      @      @      4@     �I@     �B@      B@     �B@     �A@      @@       @      $@     �@@      6@      6@      4@      4@      $@      .@      @      @      @      $@              @      @       @      $@      �?      @      �?      @      &@       @      @       @       @              �?      @      .@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ,�hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKqhth)h,K ��h.��R�(KKq��h{�B@         0                     @\H�l�?�           @�@       @       #                    �?d�2�,��?�            �r@    �8@                           (@���*~�?s            @f@ 5Y��  ������������������������       �                     ,@0Z��                              �?�p ��?k            �d@      @                          �G@�+e�X�?3            �R@    �M@                        `fpk@ {��e�?"            �J@    �E@                         x#J@r�q��?             H@       	       
                 �T!@@ �Cc}�?             <@        ������������������������       ��z�G��?	             $@      @������������������������       �        	             2@      ;@                        Ј@S@      �?             4@      �?������������������������       ����Q��?             @�                               �y[@�r����?             .@      �?������������������������       �                      @      �?������������������������       �����X�?             @      @������������������������       ����Q��?             @Z                              �D8H@�X����?             6@                              ���=@���Q��?	             $@       ������������������������       �z�G�z�?             @w      ������������������������       ����Q��?             @n      ������������������������       �      �?             (@�                                 �?���M�?8            @V@       ������������������������       �؇���X�?             @�                                �?@0��P�?3            �T@                                 &@��Y��]�?            �D@       ������������������������       �$�q-�?	             *@      ������������������������       �                     <@                                @A@������?            �D@       ������������������������       ��z�G��?             $@(             "                    �?�g�y��?             ?@              !                 ��Y)@�}�+r��?
             3@       ������������������������       �؇���X�?             @3      ������������������������       �                     (@A      ������������������������       �                     (@�       $       -                  "�b@0 �����?J            @^@       %       (                   �;@����w�?A            @[@        &       '                    6@�#-���?            �A@        ������������������������       �      �?              @�       ������������������������       �                     ;@�       )       ,                    �?`׀�:M�?*            �R@        *       +                 hf(P@�X�<ݺ?
             2@        ������������������������       �z�G�z�?             @$       ������������������������       �                     *@       ������������������������       �                      L@       .       /                 `D�g@�q�q�?	             (@        ������������������������       ��q�q�?             @]       ������������������������       �                     @�       1       >                    �?��i��?           �y@        2       9                    �?(옄��?             G@       3       4                 ���@�n_Y�K�?             :@        ������������������������       �                     @�       5       6                    ;@�\��N��?             3@        ������������������������       ������H�?             "@      7       8                   @@z�G�z�?
             $@        ������������������������       �z�G�z�?             @`      ������������������������       �z�G�z�?             @:      :       =                 ���.@      �?             4@      ;       <                    �?�q�q�?             (@       ������������������������       �r�q��?             @I      ������������������������       ��q�q�?             @7      ������������������������       �                      @G       ?       D                    @>�y@��?�            �v@       @       A                     @
;&����?             7@       ������������������������       �                     @�      B       C                    @      �?	             0@       ������������������������       �                      @8       ������������������������       �      �?              @8      E       f                   �@@�4���L�?�            �u@      F       O                 ��@2ۭVJ�?�            �q@       G       L                    �?���e��?)            �P@      H       I                 ���@�?�'�@�?             C@       ������������������������       ����!pc�?             &@�       J       K                    �?�>����?             ;@       ������������������������       �8�Z$���?             *@v      ������������������������       �                     ,@�      M       N                    9@����X�?             <@       ������������������������       �z�G�z�?             $@�      ������������������������       ��q�q�?             2@�      P       e                   �>@z�z�7��?�            `k@      Q       \                   �;@ޗQ�~�?�            �i@       R       [                   �:@p��*�?F            �[@      S       Z                    �?�DÓ ��?A            @Y@      T       U                    �?�T|n�q�?5            �U@      ������������������������       ���v����?)            �P@g      V       Y                    �?�d�����?             3@       W       X                    0@�q�q�?             .@        ������������������������       �����X�?             @}       ������������������������       �                      @�       ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                     "@        ]       d                   �=@dP-���?;            �W@       ^       _                 ��) @Du9iH��?6            �U@        ������������������������       �                    �E@        `       a                    �?(L���?            �E@        ������������������������       ��q�q�?             "@        b       c                    �?l��\��?             A@       ������������������������       �@�0�!��?             1@        ������������������������       �                     1@        ������������������������       �      �?              @        ������������������������       ���S���?             .@        g       l                 `f�"@ ,��-�?#            �M@       h       k                   �C@��Y��]�?            �D@        i       j                   �A@@4և���?	             ,@       ������������������������       �                      @        ������������������������       �r�q��?             @        ������������������������       �                     ;@        m       p                 0336@r�q��?             2@       n       o                    �?�z�G��?             $@        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                      @        �t�b�@     h�h)h,K ��h.��R�(KKqKK��h\�B       �|@     �o@     �b@     �b@     �a@      C@              ,@     �a@      8@     �L@      2@      E@      &@      D@       @      9@      @      @      @      2@              .@      @       @      @      *@       @       @              @       @       @      @      .@      @      @      @      @      �?       @      @      "@      @     �T@      @      @      �?     @S@      @      D@      �?      (@      �?      <@             �B@      @      @      @      >@      �?      2@      �?      @      �?      (@              (@               @     @\@      @     @Z@      @      @@      @      @              ;@      �?     @R@      �?      1@      �?      @              *@              L@      @       @      @       @              @     Ps@      Z@      5@      9@      0@      $@      @              "@      $@      �?       @       @       @      @      �?      @      �?      @      .@      @      @      �?      @      @       @               @      r@     �S@      (@      &@              @      (@      @       @              @      @     @q@      Q@     �k@      P@     �D@      9@     �@@      @       @      @      9@       @      &@       @      ,@               @      4@       @       @      @      (@     �f@     �C@     �e@      ?@     �U@      7@     �U@      ,@      R@      ,@      M@      "@      ,@      @      $@      @       @      @       @              @              .@                      "@     �U@       @      T@      @     �E@             �B@      @      @      @      ?@      @      ,@      @      1@              @       @      @       @     �K@      @      D@      �?      *@      �?       @              @      �?      ;@              .@      @      @      @      @              �?      @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJf��'hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK	hsKOhth)h,K ��h.��R�(KKO��h{�B�         .                    �?�}���?�           @�@      @                           $@d�!��?1           �|@ , 4.],                           �;@��H�}�?             9@  be use������������������������       �                     *@>> x1 = ������������������������       �      �?             (@      �?                            �?ZدG�<�?           @{@      �?                        ��$:@l�Ӑ���?=            �U@        ������������������������       �                     @      �?	                           �?2lK����?8            @T@     @\@
                           �?r�q��?             8@     ;@                         �}S@     ��?             0@     *@������������������������       �և���X�?             @      @������������������������       ������H�?             "@�       ������������������������       �      �?              @      �?                        ��yC@��U/��?'            �L@      @                           D@l��[B��?             =@      &@������������������������       �z�G�z�?             $@Z                                �J@�����?             3@       ������������������������       �X�<ݚ�?             "@�      ������������������������       �z�G�z�?             $@w                                 �? �Cc}�?             <@       ������������������������       �        	             *@�                                 D@z�G�z�?             .@       ������������������������       ��q�q�?             @�      ������������������������       ������H�?             "@�             '                 `��+@�4�`WC�?�            �u@             &                 ��@�x{��?�            q@              !                    �?      �?8             X@                                 �:@ܷ��?��?             =@       ������������������������       �����X�?             @(                               ���@���7�?             6@       ������������������������       �                     $@J      ������������������������       ��8��8��?             (@3      "       #                   �;@�����?&            �P@       ������������������������       ������?             5@�       $       %                   �=@��<b�ƥ?             G@        ������������������������       ����7�?             6@v       ������������������������       �                     8@j       ������������������������       �nS޸��?s             f@�       (       -                 �T�I@p�|�i�?6             S@       )       *                    �? ��ʻ��?1             Q@       ������������������������       �        )             L@�       +       ,                    :@�8��8��?             (@        ������������������������       �                     @       ������������������������       �r�q��?             @       ������������������������       �      �?              @-       /       8                     @AB����?�            `o@       0       1                    @=QcG��?T            �a@        ������������������������       �      �?              @A       2       3                    6@0�!F��?P            �`@        ������������������������       ��r����?             >@�       4       5                    �?@�n���?=            �Y@       ������������������������       �        2             U@�       6       7                   �W@�}�+r��?             3@      ������������������������       �                     $@�       ������������������������       ������H�?             "@`      9       :                  s�@�eP*L��?I            �[@       ������������������������       �                     "@;      ;       L                    @l@!���?B            @Y@      <       C                 P��%@���>4��?8             U@       =       @                   �:@���Q �?            �H@       >       ?                    3@"pc�
�?             6@        ������������������������       ����Q��?             $@      ������������������������       �                     (@!      A       B                    �?|��?���?             ;@      ������������������������       �X�Cc�?	             ,@�      ������������������������       ��	j*D�?             *@8       D       E                 P��+@<=�,S��?            �A@       ������������������������       �                      @      F       G                 �?�-@|��?���?             ;@       ������������������������       �                     @,      H       I                    �?���|���?             6@       ������������������������       �                     "@�       J       K                 ���3@�n_Y�K�?
             *@        ������������������������       �      �?              @v      ������������������������       �z�G�z�?             @�      M       N                    !@�t����?
             1@       ������������������������       ��q�q�?             @�      ������������������������       �                     &@�      �t�bh�h)h,K ��h.��R�(KKOKK��h\�B�       |@     pp@     �w@     @T@      "@      0@              *@      "@      @     0w@     @P@     �M@      <@      @             �J@      <@      *@      &@      &@      @      @      @       @      �?       @      @      D@      1@      .@      ,@       @       @      *@      @      @      @       @       @      9@      @      *@              (@      @      @       @       @      �?     �s@     �B@     �m@      A@     �V@      @      :@      @      @       @      5@      �?      $@              &@      �?      P@      @      3@       @     �F@      �?      5@      �?      8@             �b@      <@     @R@      @     �P@      �?      L@              &@      �?      @              @      �?      @       @     @Q@     �f@      "@     �`@      @      @      @      `@      @      :@      �?     �Y@              U@      �?      2@              $@      �?       @      N@      I@              "@      N@     �D@     �F@     �C@      @@      1@      2@      @      @      @      (@              ,@      *@      @      "@      "@      @      *@      6@               @      *@      ,@      @               @      ,@              "@       @      @      @      @      @      �?      .@       @      @       @      &@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJy"rhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKmhth)h,K ��h.��R�(KKm��h{�B@                          Ь�#@�?a/���?�           @�@       @                           �?    ���?�             p@rrorr
                           �;@��j�o�?�            �i@ 5H��                             �?�Y����?,            �P@ ��Ձ��������������������������       ��q�q�?             @       @������������������������       ���.��?'            �N@       @                           �?PX�V|�?X            `a@      @       	                 ���@l��\��?             A@        ������������������������       �                     @      �?
                           =@�����H�?             ;@     @                         s�@�S����?             3@        ������������������������       �ףp=
�?             $@     �`@������������������������       ��<ݚ�?             "@�       ������������������������       �                      @       @                          �C@��FM ò?D            @Z@    �C@������������������������       � �\���?4            �S@        ������������������������       �                     :@                                pF @���Q��?$             I@                               P�@�����?             C@        ������������������������       �      �?              @                                ��@������?             >@        ������������������������       �     ��?	             0@                                0�w@X�Cc�?             ,@        ������������������������       �և���X�?             @        ������������������������       �����X�?             @                                `�X!@�q�q�?
             (@        ������������������������       �                     @        ������������������������       �և���X�?             @               X                  x#J@�Uo���?            �|@              A                     @�(�k�I�?�             t@                                   .@2���?}            �g@        ������������������������       �        
             *@        !       >                   @L@����*��?s             f@      "       =                    �?�����?i            �c@      #       6                    �?�\��N��?e             c@       $       '                    �?�����??            �X@        %       &                   �<@X�Cc�?	             ,@        ������������������������       �և���X�?             @j       ������������������������       �؇���X�?             @�       (       -                     �?�>4և��?6             U@        )       ,                   �H@��
ц��?             :@       *       +                   �>@j���� �?             1@        ������������������������       �      �?              @$       ������������������������       �                     "@       ������������������������       �X�<ݚ�?             "@       .       5                    �?�8���?&             M@       /       0                    &@ "��u�?              I@        ������������������������       �z�G�z�?             $@�       1       2                   �@@�(\����?             D@       ������������������������       �                     6@�       3       4                   �B@�X�<ݺ?             2@        ������������������������       �r�q��?             @�       ������������������������       �                     (@�       ������������������������       �                      @      7       <                    �? 7���B�?&             K@       8       ;                    �?���N8�?             E@      9       :                    �?Pa�	�?            �@@       ������������������������       ��C��2(�?             &@;      ������������������������       �                     6@?      ������������������������       ������H�?             "@I      ������������������������       �        	             (@7      ������������������������       �                     @G       ?       @                     �?�����H�?
             2@      ������������������������       ��8��8��?             (@!      ������������������������       �r�q��?             @�      B       M                    �?FVQ&�?O            �`@      C       H                    *@�MI8d�?+            �R@        D       E                    @�eP*L��?             6@       ������������������������       �r�q��?             @      F       G                   X1@     ��?	             0@       ������������������������       �                     "@,      ������������������������       �                     @�      I       L                    �? ��WV�?             J@        J       K                 ��$1@8�Z$���?	             *@       ������������������������       �                      @v      ������������������������       ����Q��?             @�      ������������������������       �                    �C@�      N       O                    �?��o	��?$             M@       ������������������������       �                     @�      P       W                 ��Y7@�F�j��?             �J@      Q       T                    �?��Q��?             D@       R       S                    5@���Q��?             9@       ������������������������       �z�G�z�?             $@-      ������������������������       ��r����?	             .@%      U       V                    �?������?
             .@       ������������������������       �z�G�z�?             @�       ������������������������       ��z�G��?             $@y       ������������������������       �        	             *@}       Y       l                    @�iޤ��?T            �`@       Z       ]                    4@@�j���?N            @_@        [       \                    �?��
ц��?
             *@        ������������������������       �r�q��?             @        ������������������������       �����X�?             @        ^       i                    �?����1�?D             \@        _       h                    �?      �?             H@       `       c                    �?�G��l��?             E@        a       b                  �}S@�eP*L��?
             6@       ������������������������       �����X�?             ,@        ������������������������       �      �?              @        d       g                    �?      �?             4@       e       f                 ЈrS@���|���?
             &@        ������������������������       �      �?             @        ������������������������       �z�G�z�?             @        ������������������������       ��q�q�?             "@        ������������������������       ��q�q�?             @        j       k                    �?     ��?'             P@       ������������������������       �                    �I@        ������������������������       �$�q-�?             *@        ������������������������       �                     "@        �t�bh�h)h,K ��h.��R�(KKmKK��h\�B�        {@     �q@     �i@     �H@     `g@      3@     �K@      (@      @       @     �I@      $@     �`@      @      ?@      @      @              8@      @      0@      @      "@      �?      @       @       @             @Y@      @     �R@      @      :@              4@      >@      (@      :@      @      @       @      6@      @      *@      @      "@      @      @       @      @       @      @      @              @      @      l@     �l@      g@      a@      X@     �W@              *@      X@     @T@      T@     �S@      T@      R@     �S@      4@      "@      @      @      @      @      �?     @Q@      .@      ,@      (@      $@      @      �?      @      "@              @      @     �K@      @     �G@      @       @       @     �C@      �?      6@              1@      �?      @      �?      (@               @               @      J@       @      D@      �?      @@      �?      $@              6@      �?       @              (@              @      0@       @      &@      �?      @      �?     @V@     �E@      O@      (@      (@      $@      @      �?      @      "@              "@      @              I@       @      &@       @       @              @       @     �C@              ;@      ?@              @      ;@      :@      ,@      :@      $@      .@       @       @       @      *@      @      &@      �?      @      @      @      *@              D@     �W@      ?@     �W@      @      @      �?      @      @       @      9@     �U@      8@      8@      4@      6@      $@      (@      @      $@      @       @      $@      $@      @      @      @      @      @      �?      @      @      @       @      �?     �O@             �I@      �?      (@      "@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�A�'hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKwhth)h,K ��h.��R�(KKw��h{�B�         N                    �?<��z��?�           @�@      @                           @Ԛ��]m�?           |@ �^��                          @3�4@�t����?             1@ �e��  ������������������������       �                     "@tL�K<׮t������������������������       �      �?              @      @       A                 `fFJ@�_p�<�?            {@     @       6                   @@@     |�?�             x@     @       5                   �?@ 4�"=[�?�            �n@     *@	       
                    *@��g�g�?�            �m@      4@������������������������       �      �?              @      .@                          �8@h�˹�?�            �l@                                   �?���N8�?3             U@       @������������������������       �8�Z$���?             *@�                                 �4@�J�T�?.            �Q@     D@                           �?�7��?            �C@      @                            @��?^�k�?            �A@      �?������������������������       �                      @Z                                �2@ 7���B�?             ;@       ������������������������       �                     $@�                                �3@�IєX�?	             1@      ������������������������       �؇���X�?             @n      ������������������������       �                     $@�      ������������������������       �      �?             @�      ������������������������       �                     @@�             "                    �?�E���-�?_             b@              !                 м;4@H�ՠ&��?"             K@                                  �?���V��?            �F@                                 �?��G���?            �B@                                 @@      �?             4@      ������������������������       �"pc�
�?             &@(      ������������������������       ��q�q�?             "@V      ������������������������       ��t����?             1@J      ������������������������       �                      @3      ������������������������       �                     "@A      #       $                 `f�@:	��ʵ�?=            �V@        ������������������������       �                     "@�       %       &                   �9@|��"J�?8            @T@        ������������������������       �X�<ݚ�?             "@j       '       ,                 ��) @r�q��?4             R@        (       )                  sW@l��\��?             A@        ������������������������       ��q�q�?             @�       *       +                 @3�@h�����?             <@       ������������������������       �$�q-�?             *@$       ������������������������       �        
             .@       -       4                    �?�I�w�"�?             C@       .       3                     @8^s]e�?             =@       /       2                   �<@�<ݚ�?             2@       0       1                 `f�<@�q�q�?             (@        ������������������������       �z�G�z�?             @A       ������������������������       �և���X�?             @�       ������������������������       �                     @�       ������������������������       ��eP*L��?             &@�       ������������������������       �                     "@�       ������������������������       ��z�G��?             $@      7       >                 ��D:@p��%���?N            @a@       8       =                   �N@�|1)�?=            �Z@      9       <                    A@�eGk�T�?9            �W@       :       ;                     @�nkK�?             7@       ������������������������       �      �?              @?      ������������������������       �                     .@I      ������������������������       �        -             R@7      ������������������������       �"pc�
�?             &@G       ?       @                   �C@     ��?             @@       ������������������������       ��q�q�?             @!      ������������������������       �ȵHPS!�?             :@�      B       C                 `�jM@�q�q�?!             H@       ������������������������       ��n_Y�K�?             *@8       D       I                 03�U@4�2%ޑ�?            �A@      E       H                     �?�����?             5@      F       G                 `f�S@�r����?	             .@       ������������������������       �r�q��?             @,      ������������������������       ������H�?             "@�      ������������������������       �                     @�       J       M                    �?և���X�?             ,@       K       L                  "&d@�<ݚ�?             "@       ������������������������       �z�G�z�?             @�      ������������������������       �      �?             @�      ������������������������       �z�G�z�?             @�      O       `                     @T�MB��?�            pp@      P       ]                 ���a@`Ӹ����?Z            �`@      Q       Z                   �H@0x�!���?M            �]@       R       Y                    6@p���?D             Y@       S       X                 ��[,@�>����?             ;@      T       U                    �?���N8�?             5@       ������������������������       �                     @g      V       W                   @>@��S�ۿ?
             .@        ������������������������       �؇���X�?             @y       ������������������������       �                      @}       ������������������������       �r�q��?             @�       ������������������������       �        2            @R@        [       \                   @I@�KM�]�?	             3@        ������������������������       �      �?              @        ������������������������       �                     &@        ^       _                    �?      �?             0@       ������������������������       �                     "@        ������������������������       �����X�?             @        a       v                 ��Y7@     ^�?L             `@       b       g                 ��@�	��)��??            �Y@        c       f                 ���@��<b���?             7@       d       e                    �?؇���X�?
             ,@       ������������������������       �����X�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             "@        h       k                    �?R�����?0             T@        i       j                 03�-@�q�q�?             8@        ������������������������       ��<ݚ�?             "@        ������������������������       �        
             .@        l       q                  �#@X�Cc�?!             L@        m       p                    �?�q�q�?             8@       n       o                   �9@     ��?
             0@        ������������������������       ��<ݚ�?             "@        ������������������������       �և���X�?             @        ������������������������       �                      @        r       u                 ��1@     ��?             @@       s       t                    �?z�G�z�?             .@        ������������������������       �r�q��?             @        ������������������������       ��<ݚ�?             "@        ������������������������       �@�0�!��?             1@        ������������������������       �                     9@        �t�bh�h)h,K ��h.��R�(KKwKK��h\�Bp       p|@     p@     �w@     @R@      @      (@              "@      @      @     0w@     �N@     0u@     �F@      j@     �B@     �i@      >@      @      @      i@      ;@      T@      @      &@       @     @Q@       @     �B@       @      A@      �?       @              :@      �?      $@              0@      �?      @      �?      $@              @      �?      @@             @^@      7@     �G@      @      C@      @      >@      @      .@      @      "@       @      @      @      .@       @       @              "@             �R@      0@      "@             @P@      0@      @      @      N@      (@      ?@      @      @       @      ;@      �?      (@      �?      .@              =@      "@      4@      "@      ,@      @       @      @      @      �?      @      @      @              @      @      "@              @      @     @`@       @     �Y@      @     �W@      �?      6@      �?      @      �?      .@              R@              "@       @      ;@      @      @       @      7@      @      @@      0@      @       @      ;@       @      3@       @      *@       @      @      �?       @      �?      @               @      @      @       @      @      �?      @      �?      �?      @     �S@      g@      @      `@      @     �\@       @     �X@       @      9@      �?      4@              @      �?      ,@      �?      @               @      �?      @             @R@       @      1@       @      @              &@       @      ,@              "@       @      @     @R@     �K@      H@     �K@      @      2@       @      (@       @      @              @      @      @     �E@     �B@      @      1@      @       @              .@      B@      4@      3@      @      &@      @      @       @      @      @       @              1@      .@      @      (@      �?      @       @      @      ,@      @      9@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ���hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKchth)h,K ��h.��R�(KKc��h{�B�                             @T�����?�           @�@       @                        �Q��?p9W��S�?             C@ ���  ������������������������       �                     $@pZ8��                             @��>4և�?             <@o�4                               @�t����?             1@     �?������������������������       ��<ݚ�?             "@        ������������������������       �                      @      @������������������������       �"pc�
�?             &@       @	       <                    �?�oMo��?�           �@       
       -                  I>@�S����?           P{@     @                         s�@�Jx��?�            0v@                                ���@�&=�w��?'            �J@      @������������������������       �                     4@�                                 �;@�FVQ&�?            �@@      @������������������������       �z�G�z�?             $@        ������������������������       �                     7@       @       ,                    �?�npº��?�            �r@                                  �? B�*]-�?�            �q@                               ��";@      �?             <@      ������������������������       ��q�q�?             2@w      ������������������������       �ףp=
�?             $@n             +                 �y�/@L紂P�?�            �o@             *                    �?v&�����?�            �j@                              �1@�0]�I�?~            �i@                                  >@�E��ӭ�?             B@                                �8@�q�q�?             >@       ������������������������       �ףp=
�?             $@      ������������������������       ��G�z��?             4@      ������������������������       �                     @�                              �?�@x-B�?i             e@       ������������������������       �                    �E@V              !                 @3�@�nN@��?P            �_@       ������������������������       ��<ݚ�?             "@3      "       #                 ��i @�����8�?J            @]@       ������������������������       ��������?             F@�       $       %                 ���$@����1�?2            @R@        ������������������������       �                     ;@v       &       '                    5@*
;&���?              G@        ������������������������       �      �?             @�       (       )                    �?ףp=
�?             D@        ������������������������       �                      @�       ������������������������       �      �?             @@�       ������������������������       �����X�?             @$       ������������������������       �                    �E@       ������������������������       �        	             3@       .       7                    �?��p �?6            �T@       /       2                   �;@և���X�?!            �H@        0       1                   �9@�q�q�?	             (@       ������������������������       �և���X�?             @A       ������������������������       �                     @�       3       6                 Ј�T@^H���+�?            �B@       4       5                    �?:ɨ��?            �@@       ������������������������       ��q�q�?             8@�       ������������������������       �                     "@      ������������������������       �      �?             @�       8       9                    �?<���D�?            �@@       ������������������������       ��z�G��?             $@:      :       ;                    �?�nkK�?             7@       ������������������������       �r�q��?             @?      ������������������������       �        	             1@I      =       >                    (@�2��?�            �m@       ������������������������       ��C��2(�?             &@G       ?       L                     @
�ۓQ{�?�            @l@      @       G                 03[=@`�c�г?R             _@       A       B                    �?���}<S�?!             G@       ������������������������       �����X�?             @�      C       F                    6@�7��?            �C@       D       E                   �;@���}<S�?             7@       ������������������������       �      �?              @      ������������������������       �                     .@-      ������������������������       �                     0@,      H       I                 ���a@�(�Tw�?1            �S@      ������������������������       �        $            �N@�       J       K                    �?�IєX�?             1@       ������������������������       �                     &@v      ������������������������       �r�q��?             @�      M       `                   @B@�ʻ����?B            �Y@      N       _                    �?������?:            �U@      O       V                    �?�O�y���?3            �R@       P       S                 Ь* @�(�Tw��?            �C@      Q       R                   �2@�LQ�1	�?             7@        ������������������������       �                     @      ������������������������       ��S����?
             3@-      T       U                 ��.@      �?	             0@      ������������������������       �                      @g      ������������������������       �                      @�       W       ^                   �>@*O���?             B@       X       [                   �;@¦	^_�?             ?@       Y       Z                  �#@j���� �?             1@       ������������������������       ��z�G��?             $@        ������������������������       �և���X�?             @        \       ]                    �?؇���X�?
             ,@        ������������������������       �                     @        ������������������������       �����X�?             @        ������������������������       �z�G�z�?             @        ������������������������       �r�q��?             (@        a       b                    E@�r����?             .@        ������������������������       �                     "@        ������������������������       ��q�q�?             @        �t�bh�h)h,K ��h.��R�(KKcKK��h\�B0       0|@     Pp@      &@      ;@              $@      &@      1@       @      .@       @      @               @      "@       @     �{@     @m@      w@     @Q@     ps@      F@     �I@       @      4@              ?@       @       @       @      7@             @p@      E@      n@      E@      5@      @      (@      @      "@      �?     �k@     �A@      f@     �A@     �e@     �@@      :@      $@      4@      $@      "@      �?      &@      "@      @             @b@      7@     �E@             �Y@      7@       @      @     @Y@      0@     �A@      "@     �P@      @      ;@             �C@      @      @      @      B@      @       @              <@      @      @       @     �E@              3@             �L@      9@      <@      5@      @       @      @      @              @      8@      *@      7@      $@      ,@      $@      "@              �?      @      =@      @      @      @      6@      �?      @      �?      1@              R@     �d@      $@      �?      O@     �d@      @     �]@      @      E@       @      @       @     �B@       @      5@       @      @              .@              0@      �?     @S@             �N@      �?      0@              &@      �?      @     �L@     �F@      F@     �E@      A@     �D@      &@      <@      @      4@              @      @      0@       @       @       @                       @      7@      *@      6@      "@      $@      @      @      @      @      @      (@       @      @              @       @      �?      @      $@       @      *@       @      "@              @       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJJ��hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKhth)h,K ��h.��R�(KK��h{�B�         8                     @�)�>_M�?�           @�@       @                           �?և���X�?�            �r@ �Ġ�                             �?���5��?0            �S@1���                             �?$]��<C�?+            �Q@ 2���                          �ܵ<@���@M^�?             ?@        ������������������������       �                     @               
                    �?l��
I��?             ;@              	                 `f�B@�q�q�?
             5@        ������������������������       �z�G�z�?             .@        ������������������������       ��q�q�?             @        ������������������������       �r�q��?             @                                ��A@P���Q�?             D@        ������������������������       �      �?              @        ������������������������       �                     @@        ������������������������       �և���X�?             @                                  �.@�[����?�            �k@                                   �?r֛w���?+             O@{���s�                           &@�t����?#            �I@ n���9                           @������?             1@�q��r=�������������������������       �                     "@���W�b9������������������������       �      �?              @ gL��g*(                        `f�)@�IєX�?             A@ G͊����������������������������       �                     @w�Q��                           =@�>����?             ;@ '�l�Y�                          �8@؇���X�?	             ,@ ԥ>��eK������������������������       �                     @T�#M����������������������������       ��<ݚ�?             "@��[�D�������������������������       �        	             *@m�~����                           :@�C��2(�?             &@ ���AY��������������������������       �z�G�z�?             @@>7]�hn������������������������       �                     @��V�נ�        1                    �?ZSu6��?g             d@Y�}�0ԩ!       0                  D0T@�A����?8            �T@      "       #                    %@^��4m�?3            �R@       ������������������������       �                     @�       $       -                   @E@�Y����?/            �P@       %       &                 ��D:@�θ�?            �C@        ������������������������       �                     $@j       '       ,                     �?8^s]e�?             =@       (       +                   �@@և���X�?             5@       )       *                 �T9G@������?             .@        ������������������������       ��q�q�?             @�       ������������������������       ��<ݚ�?             "@$       ������������������������       �r�q��?             @       ������������������������       �                      @       .       /                   �G@ �Cc}�?             <@        ������������������������       �                     $@]       ������������������������       �r�q��?             2@�       ������������������������       �      �?              @A       2       7                   �;@p`q�q��?/            �S@        3       4                     �?�'�`d�?            �@@        ������������������������       ���
ц��?             *@�       5       6                    :@P���Q�?             4@        ������������������������       �ףp=
�?             $@      ������������������������       �                     $@�       ������������������������       �                     G@`      9       `                    �?�:���?           �y@      :       _                 �T�I@�ˡ�5��?�            �q@      ;       \                    @8�Z$���?�            q@      <       =                   �0@    �7�?�             p@       ������������������������       ��q�q�?             (@7      >       W                   @@@��̋���?�            �n@       ?       D                 �Y�@�s�;�w�?w            �f@       @       C                    �?����X�?            �A@      A       B                 ���@�����?             3@       ������������������������       �؇���X�?             @�      ������������������������       ��q�q�?             (@8       ������������������������       �      �?             0@8      E       F                    �?�x
�2�?d            �b@       ������������������������       �z�G�z�?             $@-      G       L                   �:@�θV�?`            @a@       H       K                   �4@�1�`jg�?$            �K@       I       J                 P�@�S����?             3@        ������������������������       �                     "@�       ������������������������       ��z�G��?             $@v      ������������������������       �                     B@�      M       R                   �@�o��gn�?<            �T@       N       Q                 ��@d}h���?             <@      O       P                 03�@�C��2(�?             6@       ������������������������       �                     $@�      ������������������������       �r�q��?             (@�       ������������������������       ��q�q�?             @      S       V                    �?�C��2(�?+            �K@      T       U                   �>@ףp=
�?!             D@      ������������������������       ��FVQ&�?            �@@g      ������������������������       �����X�?             @�       ������������������������       ���S�ۿ?
             .@y       X       Y                   �E@�]0��<�?&            �N@       ������������������������       �                    �D@�       Z       [                   �G@ףp=
�?             4@        ������������������������       �      �?              @        ������������������������       �        	             (@        ]       ^                    �?�IєX�?             1@       ������������������������       �                     &@        ������������������������       �r�q��?             @        ������������������������       ��eP*L��?             &@        a       l                    �?b7s�H�?R            �_@        b       e                   �0@���Q��?             I@        c       d                   �+@�8��8��?             (@        ������������������������       �                     @        ������������������������       �r�q��?             @        f       k                 ��.@      �?             C@       g       h                    9@     ��?             @@        ������������������������       ��q�q�?             "@        i       j                    �?\X��t�?             7@        ������������������������       ��q�q�?             @        ������������������������       ���.k���?
             1@        ������������������������       �                     @        m       v                   �7@��cv�?4            @S@        n       q                    �?և���X�?            �A@        o       p                 �&B@p�ݯ��?             3@        ������������������������       �                     "@        ������������������������       ��z�G��?             $@        r       u                    ,@     ��?             0@       s       t                    @ףp=
�?	             $@       ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       ��q�q�?             @        w       |                   �>@d}h���?             E@       x       y                   �&@��� ��?             ?@        ������������������������       �                     *@        z       {                 pf�2@�<ݚ�?             2@        ������������������������       ��q�q�?             @        ������������������������       �                     (@        }       ~                   �C@�eP*L��?             &@        ������������������������       �r�q��?             @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KKKK��h\�B�       `{@      q@      `@     �e@      1@     �N@      ,@     �L@      (@      3@      @               @      3@      @      ,@      @      (@      @       @      �?      @       @      C@       @      @              @@      @      @      \@     �[@      G@      0@     �F@      @      *@      @      "@              @      @      @@       @      @              9@       @      (@       @      @              @       @      *@              �?      $@      �?      @              @     �P@     �W@     �M@      7@     �K@      3@              @     �K@      (@      >@      "@      $@              4@      "@      (@      "@      &@      @      @       @      @       @      �?      @       @              9@      @      $@              .@      @      @      @      @      R@      @      :@      @      @      �?      3@      �?      "@              $@              G@     Ps@     �Y@     �m@      H@     �l@      E@     �j@     �D@      @      @     @j@      A@     �b@      @@      9@      $@      *@      @      @      �?      @      @      (@      @     �_@      6@       @       @      _@      ,@      J@      @      0@      @      "@              @      @      B@              R@      &@      6@      @      4@       @      $@              $@       @       @      @      I@      @      B@      @      ?@       @      @       @      ,@      �?     �M@       @     �D@              2@       @      @       @      (@              0@      �?      &@              @      �?      @      @     @R@      K@      4@      >@      �?      &@              @      �?      @      3@      3@      3@      *@      @      @      *@      $@      @       @      "@       @              @     �J@      8@      4@      .@      @      (@              "@      @      @      *@      @      "@      �?      @              @      �?      @       @     �@@      "@      ;@      @      *@              ,@      @       @      @      (@              @      @      �?      @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�U�uhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKehth)h,K ��h.��R�(KKe��h{�B@         (                     @r�����?�           @�@       @                         x#J@� �	��?�            Pt@                                  �?$_;|��?�            �j@                               ��D:@\�CX�?Y            �a@                                  �?,���i�?4            �T@       ������������������������       �@݈g>h�?0             S@        ������������������������       �      �?             @                                  �?@d��0u��?%             N@       	       
                 ���<@�������?             >@        ������������������������       �                      @                                   �?�X����?             6@       ������������������������       ��n_Y�K�?             *@        ������������������������       ��<ݚ�?             "@                                �T!@@      �?             >@                                 �J@�q�q�?             8@                                �C@      �?             0@        ������������������������       �����X�?             @Z      ������������������������       ��<ݚ�?             "@�      ������������������������       �      �?              @�      ������������������������       �r�q��?             @w                                  �?0z�(>��?+            �Q@       ������������������������       �"pc�
�?             &@�                              ���*@ �.�?Ƞ?%             N@                                  =@���7�?             6@       ������������������������       ��C��2(�?             &@�      ������������������������       �                     &@c      ������������������������       �                     C@                                �1@���X�?F             \@       ������������������������       �                     (@�             '                    �?�z�G��??             Y@                                  �8@����X�?             E@       ������������������������       �                     @J      !       "                 03�M@^������?            �A@       ������������������������       �z�G�z�?             @A      #       $                 �U�R@������?             >@        ������������������������       �                      @�       %       &                 ���X@���|���?             6@        ������������������������       ���
ц��?             *@j       ������������������������       ������H�?             "@�       ������������������������       �        "             M@�       )       L                    �?���t�?�            0x@       *       /                    *@������?�            �o@        +       ,                     @r�q��?             8@        ������������������������       ��<ݚ�?             "@       -       .                    @������?             .@        ������������������������       �      �?              @-       ������������������������       �                     @]       0       1                    �?�p����?�            �l@        ������������������������       �J�8���?             =@A       2       C                   �<@�?�߾�?�             i@       3       @                 03�6@�x�+���?_            @b@       4       5                   �0@$Q�q�?T            �_@        ������������������������       �      �?              @�       6       7                   �8@����˵�?O            �]@       ������������������������       �        !            �H@�       8       ;                   �;@���}<S�?.            @Q@       9       :                 ��L@X�Cc�?             ,@       ������������������������       �և���X�?             @;      ������������������������       �؇���X�?             @?      <       ?                 �?$@ �Jj�G�?#            �K@       =       >                    �?���7�?             6@      ������������������������       �                     .@G       ������������������������       �؇���X�?             @      ������������������������       �                    �@@!      A       B                    @R���Q�?             4@      ������������������������       ����!pc�?             &@�      ������������������������       �                     "@8       D       G                   @@@�+$�jP�?%             K@       E       F                 pff@      �?             0@       ������������������������       �      �?             @-      ������������������������       ��q�q�?             (@,      H       K                 @3�@�}�+r��?             C@      I       J                 �?�@�t����?             1@       ������������������������       �        
             *@�       ������������������������       �      �?             @v      ������������������������       �                     5@�      M       d                    @B�
k���?M            �`@      N       Q                    @��Z
H��?I            @_@       O       P                 pfV0@8�Z$���?             *@       ������������������������       ��q�q�?             @�      ������������������������       �                     @�       R       S                    (@�Cc}��?A             \@       ������������������������       �                     @-      T       W                    3@Ć��H��?=            �Z@       U       V                 @1#@p�ݯ��?             3@      ������������������������       ��θ�?             *@�       ������������������������       ��q�q�?             @y       X       c                 ��Y7@ 9�����?2             V@       Y       Z                   �5@���A��?,            �R@        ������������������������       �      �?              @        [       `                   �<@����e��?'            �P@       \       ]                 ���@�I� �?             G@        ������������������������       ��8��8��?             (@        ^       _                 pF�-@j���� �?             A@       ������������������������       �8�A�0��?             6@        ������������������������       ��8��8��?             (@        a       b                    A@�G�z��?
             4@       ������������������������       �      �?             (@        ������������������������       �      �?              @        ������������������������       �                     ,@        ������������������������       �                     "@        �t�bh�h)h,K ��h.��R�(KKeKK��h\�BP       �z@      r@     �a@     �f@     @\@      Y@     �[@      @@      R@      $@     @Q@      @      @      @      C@      6@      7@      @       @              .@      @       @      @      @       @      .@      .@      $@      ,@      @      (@       @      @       @      @      @       @      @      �?      @      Q@       @      "@      �?     �M@      �?      5@      �?      $@              &@              C@      >@     �T@              (@      >@     �Q@      >@      (@      @              7@      (@      �?      @      6@       @       @              ,@       @      @      @       @      �?              M@     �q@     �Z@     `j@      E@      *@      &@       @      @      &@      @      @      @      @             �h@      ?@      3@      $@     `f@      5@     �`@      &@     �]@       @      @       @      \@      @     �H@             �O@      @      "@      @      @      @      @      �?      K@      �?      5@      �?      .@              @      �?     �@@              1@      @       @      @      "@              F@      $@       @       @      @      �?      @      @      B@       @      .@       @      *@               @       @      5@             �Q@      P@     �N@      P@       @      &@       @      @              @     �M@     �J@      @              K@     �J@      @      (@      @      $@      @       @     �G@     �D@     �@@     �D@      @      �?      :@      D@      .@      ?@      �?      &@      ,@      4@      *@      "@      �?      &@      &@      "@      @      @      @      @      ,@              "@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJW��]hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK
hsK_hth)h,K ��h.��R�(KK_��h{�B�         <                    �?�Qc�!�?�           @�@      @       )                 ��$:@>��O�V�?*           P}@     6@       "                    �?�-q���?�            �u@     @       !                    �?��i����?�            �q@     (@                        ���#@�O��/�?�            `q@     �?                        �?�@t(d��?�            @i@     5@                          �9@4�0_���?P            @\@     �T@                          �5@�+e�X�?             9@       	       
                   �4@�8��8��?             (@       ������������������������       �                     @      M@������������������������       �z�G�z�?             @      @                          �7@�n_Y�K�?	             *@      ?@������������������������       ����Q��?             @       @������������������������       �      �?              @      @                        ���@�zvܰ?<             V@      �?������������������������       �                     F@                                   �?t��ճC�?             F@       ������������������������       ����N8�?             5@�                                �@���}<S�?             7@       ������������������������       �z�G�z�?             $@w      ������������������������       �        
             *@n      ������������������������       �&<k����?3            @V@�                                 �?p�|�i�?,             S@       ������������������������       �                     @�                                 @A@0z�(>��?(            �Q@                                  @      �?             H@                                 &@$�q-�?            �C@       ������������������������       ��C��2(�?             &@                                �;@@4և���?             <@      ������������������������       �                     4@(      ������������������������       �      �?              @V      ������������������������       �                     "@J      ������������������������       �                     7@3      ������������������������       �z�G�z�?             @A      #       $                    +@     8�?)             P@        ������������������������       �z�G�z�?             $@�       %       &                    �?�X�<ݺ?#             K@        ������������������������       �      �?              @j       '       (                 P�@�nkK�?             G@        ������������������������       ��q�q�?             @�       ������������������������       �                     D@�       *       ;                  D�\@8��~P�?N            �^@       +       6                     �?��l���?G            �[@       ,       5                    �?�����?2            �S@       -       .                   �>@\X��t�?,            @Q@        ������������������������       �*;L]n�?             >@-       /       0                 `fFJ@�q�q�?            �C@        ������������������������       ��IєX�?             1@�       1       4                   �D@�eP*L��?             6@       2       3                 `f�N@     ��?
             0@        ������������������������       �؇���X�?             @�       ������������������������       �X�<ݚ�?             "@�       ������������������������       �r�q��?             @�       ������������������������       �z�G�z�?             $@      7       :                 �T�I@�חF�P�?             ?@       8       9                    @      �?             0@       ������������������������       �r�q��?             @:      ������������������������       �                     $@;      ������������������������       �������?
             .@?      ������������������������       �r�q��?             (@I      =       H                     @ڤ���?�            `n@      >       E                    �?`���i��?T            �`@       ?       D                   �8@����X�?H             \@       @       C                    �? 7���B�?             ;@      A       B                    �?      �?
             0@       ������������������������       �                     @�      ������������������������       ������H�?             "@8       ������������������������       �        	             &@8      ������������������������       �        5            @U@      F       G                   �8@ףp=
�?             4@      ������������������������       �                     .@,      ������������������������       ����Q��?             @�      I       P                    �?��+��?C            �[@        J       K                 ���@@�0�!��?             A@        ������������������������       �                     $@v      L       O                 03�-@      �?             8@      M       N                 �&B@���Q��?             .@      ������������������������       �      �?              @�      ������������������������       �և���X�?             @�      ������������������������       �                     "@�      Q       R                 ���@�w�r��?-            @S@        ������������������������       �                     @      S       Z                    �?��M��?)            �Q@      T       Y                    �?��i#[�?             E@      U       X                   p"@�q�q�?             >@      V       W                   �9@@�0�!��?
             1@        ������������������������       �                      @y       ������������������������       ��q�q�?             "@}       ������������������������       ���
ц��?             *@�       ������������������������       �      �?             (@        [       \                 `f7@>���Rp�?             =@        ������������������������       �      �?             (@        ]       ^                    +@�IєX�?             1@        ������������������������       �      �?             @        ������������������������       �                     *@        �t�bh�h)h,K ��h.��R�(KK_KK��h\�B�       �{@     �p@     �w@     �U@     0s@      D@     �o@      =@     @o@      <@      f@      9@      Z@      "@      3@      @      &@      �?      @              @      �?       @      @      @       @      @      @     @U@      @      F@             �D@      @      4@      �?      5@       @       @       @      *@             @R@      0@     @R@      @      @              Q@      @     �F@      @      B@      @      $@      �?      :@       @      4@              @       @      "@              7@              @      �?     �J@      &@       @       @     �I@      @      @      �?      F@       @      @       @      D@             �R@     �G@     @R@     �B@     �G@      @@     �C@      >@      *@      1@      :@      *@      0@      �?      $@      (@      @      &@      �?      @      @      @      @      �?       @       @      :@      @      .@      �?      @      �?      $@              &@      @       @      $@      N@     �f@      @      `@      �?     �[@      �?      :@      �?      .@              @      �?       @              &@             @U@       @      2@              .@       @      @     �L@      K@      @      <@              $@      @      2@      @      "@       @      @      @      @              "@     �I@      :@              @     �I@      4@      =@      *@      4@      $@      ,@      @       @              @      @      @      @      "@      @      6@      @      @      @      0@      �?      @      �?      *@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJt�mUhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKohth)h,K ��h.��R�(KKo��h{�B�         P                    �?�Qc�!�?�           @�@      @                           @z�G�z�?%           `}@      �?                        @3�4@���N8�?             5@        ������������������������       �                     "@^��X�������������������������       ��q�q�?             (@       @                            �?�?�̌_�?           |@                                   �?J`mL�#�?;            @X@     �?                           �?�{ /h��?.            �S@       	                          �D@�4��?&            @P@      @
                          �<@�<ݚ�?             B@       @                        `fF:@P���Q�?             4@     @@������������������������       �                     &@      �?������������������������       ������H�?             "@      @                        `f�B@     ��?             0@      �?������������������������       �      �?              @      $@������������������������       �      �?              @      :@                          �J@l��[B��?             =@       ������������������������       �z�G�z�?             .@        ������������������������       �؇���X�?             ,@                                  �D@��
ц��?             *@        ������������������������       �      �?             @        ������������������������       �և���X�?             @                                03�R@�d�����?             3@        ������������������������       ��q�q�?             @                                  �E@�θ�?	             *@        ������������������������       ��q�q�?             @        ������������������������       �؇���X�?             @                                �� @      �?�             v@        ������������������������       �X�<ݚ�?             "@               O                 �T�I@�x=Fh_�?�            pu@              N                   @E@�*/�8V�?�            �t@               M                   @D@\���B��?�            �q@       !       L                    :@����?�            q@      "       #                 ���@�C͑V�?�            �o@       ������������������������       �        	             0@�       $       %                 �Y�@�v�t���?�            �m@        ������������������������       ������?             3@v       &       '                  s�@�Ra����?�            �k@        ������������������������       �                     9@�       (       A                   �<@�ݜ�?�            `h@       )       .                   @@�1�hP	�?d            �a@        *       -                 �?$@��<b���?             7@       +       ,                    ;@      �?             0@        ������������������������       �                     @       ������������������������       ��<ݚ�?             "@       ������������������������       �և���X�?             @-       /       @                    �?�8��8��?S             ^@       0       1                 �?�@l�b�G��?O            �\@        ������������������������       �                     ;@A       2       3                   �2@���(`�?>            �U@        ������������������������       �                     *@�       4       5                   �4@������?3            �R@        ������������������������       ����!pc�?             &@�       6       7                 ��) @�[|x��?+            �O@       ������������������������       �        	             *@�       8       9                   �9@ףp=
�?"             I@       ������������������������       �        
             ,@:      :       ?                    �?4?,R��?             B@      ;       >                 ���,@���B���?             :@      <       =                     @�	j*D�?
             *@       ������������������������       �����X�?             @7      ������������������������       ��q�q�?             @G       ������������������������       �$�q-�?             *@      ������������������������       �                     $@!      ������������������������       ��q�q�?             @�      B       G                   @@@���B���?"             J@       C       D                     @l��
I��?             ;@        ������������������������       �����X�?             @8      E       F                 @3�@�z�G��?             4@      ������������������������       �r�q��?             (@-      ������������������������       �      �?              @,      H       I                     @HP�s��?             9@       ������������������������       �؇���X�?             @�       J       K                 @3�@�X�<ݺ?             2@        ������������������������       �      �?              @v      ������������������������       �                     $@�      ������������������������       �                     2@�      ������������������������       ����|���?             &@�      ������������������������       �                    �F@�      ������������������������       �X�Cc�?	             ,@�      Q       Z                     @���!pc�?�            @n@       R       W                    �?�-�[�?R            ``@      S       V                    �?@3����?D             [@       T       U                   �E@�FVQ&�?            �@@      ������������������������       �                     ;@g      ������������������������       ��q�q�?             @�       ������������������������       �        .            �R@y       X       Y                 ���`@��+7��?             7@       ������������������������       �                     &@�       ������������������������       �      �?             (@        [       ^                    @�f��`��?H            �[@        \       ]                    �?     ��?             0@        ������������������������       �"pc�
�?             &@        ������������������������       �z�G�z�?             @        _       f                    �?D�n�3�?@            �W@        `       e                 ��.@�<ݚ�?             B@       a       d                 �{&@����X�?             <@       b       c                    1@"pc�
�?             6@        ������������������������       �                     @        ������������������������       �������?             .@        ������������������������       ��q�q�?             @        ������������������������       �                      @        g       j                    �?$gv&��?'            �M@        h       i                 `��!@���Q��?             4@       ������������������������       ����Q��?             $@        ������������������������       �z�G�z�?             $@        k       n                 ���4@��-�=��?            �C@        l       m                 ��Y.@���y4F�?             3@        ������������������������       �                     $@        ������������������������       �X�<ݚ�?             "@        ������������������������       �                     4@        �t�b��     h�h)h,K ��h.��R�(KKoKK��h\�B�       �{@     �p@     �w@     �W@      @      0@              "@      @      @     0w@     �S@     �O@      A@     �H@      =@     �E@      6@      <@       @      3@      �?      &@               @      �?      "@      @       @      @      @      �?      .@      ,@      @      (@      (@       @      @      @      @      @      @      @      ,@      @      @       @      $@      @      @       @      @      �?     @s@      F@      @      @     �r@      D@     `r@     �A@      o@     �A@     @n@      ?@      l@      ?@      0@              j@      ?@      *@      @     `h@      9@      9@             @e@      9@      `@      .@      2@      @      ,@       @      @              @       @      @      @     �[@      $@     �Z@       @      ;@             �S@       @      *@             �P@       @       @      @      M@      @      *@             �F@      @      ,@              ?@      @      5@      @      "@      @      @       @      @       @      (@      �?      $@              @       @      E@      $@      3@       @      @       @      ,@      @      $@       @      @      @      7@       @      @      �?      1@      �?      @      �?      $@              2@              @      @     �F@              "@      @     �P@      f@       @     �^@       @     �Z@       @      ?@              ;@       @      @             �R@      @      1@              &@      @      @      M@     �J@      @      *@       @      "@      �?      @     �K@      D@       @      <@       @      4@      @      2@              @      @      &@      @       @               @     �G@      (@      (@       @      @      @       @       @     �A@      @      .@      @      $@              @      @      4@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJc��hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKshth)h,K ��h.��R�(KKs��h{�B�         P                    �?�uY0�l�?�           @�@      @                           �?(�
��H�?.           �~@                                  �:@�J�T�?-            �Q@                                   �?և���X�?             5@                                 �6@      �?	             0@     @������������������������       �      �?              @       @������������������������       �      �?              @      F@������������������������       �z�G�z�?             @     �A@	                        ��L@@H.�!���?             I@     ?@
                            @<���D�?            �@@      9@������������������������       �8�Z$���?             *@                                  @<@ףp=
�?             4@      @������������������������       �8�Z$���?	             *@       @������������������������       �                     @      @                        ��+T@j���� �?             1@      @������������������������       �      �?             @        ������������������������       ��	j*D�?             *@Z                                 �?Dߜ���?           z@                                  �?`Ql�R�?            �G@      ������������������������       �h�����?             <@w      ������������������������       �        
             3@n                                 �?P�(ڲi�?�             w@       ������������������������       �r�q��?             @�             O                   �N@Ĝ�oV4�?�            �v@             N                  D0T@�+I�9��?�            @v@             K                    �?��	= ��?�            �u@             "                     �?ܷ��?��?�            �s@              !                 03�M@���V��?            �F@                                 @C@��G���?            �B@                                �<@����X�?             5@      ������������������������       �������?             .@V      ������������������������       ��q�q�?             @J      ������������������������       �      �?
             0@3      ������������������������       �                      @A      #       H                    �?���	���?�             q@       $       3                     @��-���?�            @p@        %       2                   �E@HP�s��?*            �R@       &       1                    �?\#r��?"            �N@       '       .                    @@$�q-�?             J@       (       )                    5@�X�<ݺ?             B@        ������������������������       �      �?              @�       *       +                   �;@h�����?             <@        ������������������������       �                     ,@$       ,       -                   �'@@4և���?             ,@        ������������������������       �                      @       ������������������������       �r�q��?             @-       /       0                   �A@      �?	             0@        ������������������������       �r�q��?             @�       ������������������������       �ףp=
�?             $@A       ������������������������       ��<ݚ�?             "@�       ������������������������       �                     ,@�       4       G                   @@@(L�\�?r             g@       5       F                    �?ϲ���?Z            �a@       6       E                   P3@��5QaJ�?R             `@      7       8                 ���@����X��?N            �^@        ������������������������       �����X�?             ,@`      9       D                   �?@|�n��T�?G            @[@      :       =                 �1@X�?٥�?C            �Y@       ;       <                 �?$@      �?             8@      ������������������������       �                     3@I      ������������������������       ����Q��?             @7      >       ?                 @3�@pY���D�?4            �S@        ������������������������       �                     <@      @       C                   �<@`'�J�?"            �I@      A       B                   �1@��<b�ƥ?             G@       ������������������������       �؇���X�?             @�      ������������������������       �                    �C@8       ������������������������       �z�G�z�?             @8      ������������������������       �r�q��?             @      ������������������������       �      �?             @-      ������������������������       �                     *@,      ������������������������       �                    �E@�      I       J                    �?d}h���?
             ,@       ������������������������       �      �?              @�       ������������������������       �                     @v      L       M                    �? 7���B�?             ;@      ������������������������       �        	             1@�      ������������������������       �ףp=
�?             $@�      ������������������������       ����Q��?             $@�      ������������������������       �      �?              @�      Q       ^                     @���X�?�             l@       R       [                   �H@P���Q�?O             ^@      S       Z                   �;@ 7���B�?F             [@       T       Y                   �8@������?            �B@      U       V                    -@��S�ۿ?             >@       ������������������������       �z�G�z�?             @�       W       X                     �?`2U0*��?             9@       ������������������������       �                     2@}       ������������������������       �؇���X�?             @�       ������������������������       �����X�?             @        ������������������������       �        ,            �Q@        \       ]                 83F@r�q��?	             (@        ������������������������       ����Q��?             @        ������������������������       �                     @        _       `                    �?��B����?H             Z@        ������������������������       �      �?             @@        a       n                    �?*O���?3             R@       b       m                   �>@X�<ݚ�?%             K@       c       h                    �?�G�z�?             D@        d       g                 ��L$@      �?             4@       e       f                 P�@�	j*D�?
             *@        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �؇���X�?             @        i       j                   @.@R���Q�?             4@        ������������������������       �                      @        k       l                    �?      �?	             (@       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �d}h���?	             ,@        o       p                    �?�����H�?             2@        ������������������������       �r�q��?             @        q       r                    +@�8��8��?             (@        ������������������������       �                      @        ������������������������       �      �?             @        �t�bh�h)h,K ��h.��R�(KKsKK��h\�B0       �}@     �m@     �y@     @R@      H@      7@      "@      (@       @       @      @      @      @      @      �?      @     �C@      &@      =@      @      &@       @      2@       @      &@       @      @              $@      @      �?      @      "@      @     �v@      I@      G@      �?      ;@      �?      3@             t@     �H@      �?      @      t@      F@     �s@      D@     �s@      A@     �q@     �@@      C@      @      >@      @      .@      @      &@      @      @       @      .@      �?       @              o@      :@     �m@      7@     @Q@      @     �K@      @      H@      @      A@       @      @      �?      ;@      �?      ,@              *@      �?       @              @      �?      ,@       @      @      �?      "@      �?      @       @      ,@              e@      1@     @_@      1@      \@      1@     @[@      ,@      $@      @     �X@      $@     �X@      @      5@      @      3@               @      @     @S@       @      <@             �H@       @     �F@      �?      @      �?     �C@              @      �?      �?      @      @      @      *@             �E@              &@      @      @      @      @              :@      �?      1@              "@      �?      @      @      @      @      N@     �d@      @     �\@      @      Z@      @     �@@       @      <@      �?      @      �?      8@              2@      �?      @       @      @             �Q@       @      $@       @      @              @      K@      I@       @      8@      G@      :@      >@      8@      ;@      *@      $@      $@      "@      @       @      @      @              �?      @      1@      @       @              "@      @      @      @      @              @      &@      0@       @      @      �?      &@      �?       @              @      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJg�$hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKqhth)h,K ��h.��R�(KKq��h{�B@         H                    �?(����7�?�           @�@      @                           �?�܆!�t�?"           �|@      �?                        xCQ@�ģ�a@�?0            @U@Q2	�                             ;@�̚��?&            �N@ �|��                             +@������?             1@      �?������������������������       �؇���X�?             @      F@������������������������       ��z�G��?             $@      @       	                     �?�Ra����?             F@       @������������������������       �������?             .@      7@
                          @@XB���?             =@      @������������������������       �                     2@      �?������������������������       ��C��2(�?             &@      �?                          �D@      �?
             8@      1@������������������������       �@�0�!��?             1@      @������������������������       �և���X�?             @                                   $@�r����?�            pw@       @                        @3�4@      �?             0@       ������������������������       �                     @�      ������������������������       ��q�q�?             "@�             ;                 `ff:@�c-vX�?�            pv@             :                    �?��� =�?�             q@                                 �?`X�Ɓ5�?�            p@       ������������������������       �XB���?             =@�             3                    &@x�}b~|�?�            �l@             2                    �?���C��?l            �c@                                  �?�KM�]�?f             c@       ������������������������       �                     @             !                   �3@L������?b            @b@                                  �2@      �?             8@                              ��Y @؇���X�?	             ,@      ������������������������       �����X�?             @V      ������������������������       �                     @J      ������������������������       ����Q��?             $@3      "       #                   �8@85�}C�?S            �^@       ������������������������       �                     ;@�       $       )                   �@�KM�]�?B            �W@        %       &                   �;@д>��C�?             =@        ������������������������       ����Q��?             @j       '       (                 P��@�8��8��?             8@       ������������������������       �                     3@�       ������������������������       ����Q��?             @�       *       /                   �?@�U�=���?+            �P@       +       .                   �<@ףp=
�?             D@       ,       -                 ��) @�IєX�?             A@       ������������������������       �                     :@       ������������������������       �      �?              @-       ������������������������       ��q�q�?             @]       0       1                 @3�@ ��WV�?             :@        ������������������������       �؇���X�?             @A       ������������������������       �                     3@�       ������������������������       �����X�?             @�       4       9                 039@��.N"Ҭ?-            @Q@       5       8                    =@P����?&            �M@       6       7                   �+@(;L]n�?             >@      ������������������������       ���S�ۿ?             .@�       ������������������������       �        
             .@`      ������������������������       �                     =@:      ������������������������       �ףp=
�?             $@;      ������������������������       �        
             .@?      <       C                    �?&[i`��?2            �U@      =       B                     @�q�q�?             H@      >       A                   �>@      �?             D@        ?       @                   �I@�\��N��?
             3@      ������������������������       ��	j*D�?             *@!      ������������������������       �r�q��?             @�      ������������������������       �                     5@�      ������������������������       �      �?              @8       D       E                   @B@$�q-�?            �C@      ������������������������       �                     9@      F       G                    �?d}h���?	             ,@      ������������������������       �����X�?             @,      ������������������������       �؇���X�?             @�      I       p                    @0,Tg��?�            �o@       J       c                 Ь�9@���?�            �n@       K       N                     @�T��5m�?O            �`@       L       M                    �?��S�ۿ?             >@      ������������������������       � ��WV�?             :@�      ������������������������       �      �?             @�      O       X                    �?��WV��?:             Z@       P       W                 ��.@�t����?            �I@      Q       V                 P��+@��]�T��?            �D@       R       S                 ��@������?             A@       ������������������������       �X�<ݚ�?             "@-      T       U                    9@�J�4�?             9@       ������������������������       �؇���X�?             @g      ������������������������       �r�q��?	             2@�       ������������������������       �                     @y       ������������������������       �                     $@}       Y       ^                   �;@l`N���?            �J@       Z       [                 pf� @�5��?             ;@        ������������������������       ����!pc�?             &@        \       ]                    �?      �?
             0@        ������������������������       �����X�?             @        ������������������������       ��q�q�?             "@        _       `                   �&@�θ�?             :@        ������������������������       �$�q-�?             *@        a       b                 03c4@�n_Y�K�?	             *@       ������������������������       �X�<ݚ�?             "@        ������������������������       �      �?             @        d       i                    �? �Cc}�?J             \@       e       h                 03[=@�e���@�?5            @S@        f       g                     �?�}�+r��?             3@        ������������������������       �r�q��?             @        ������������������������       �                     *@        ������������������������       �        )             M@        j       m                    �?">�֕�?            �A@       k       l                     �?P���Q�?             4@        ������������������������       �r�q��?             @        ������������������������       �        	             ,@        n       o                   �2@�q�q�?             .@        ������������������������       �      �?              @        ������������������������       �����X�?             @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KKqKK��h\�B       �{@      q@     `w@     �U@     �H@      B@     �E@      2@      @      *@      �?      @      @      @     �C@      @      &@      @      <@      �?      2@              $@      �?      @      2@      @      ,@      @      @     Pt@      I@      @      $@              @      @      @     �s@      D@     `o@      5@     �m@      5@      <@      �?      j@      4@     �a@      2@      a@      0@      @             @`@      0@      2@      @      (@       @      @       @      @              @      @      \@      $@      ;@             @U@      $@      8@      @       @      @      6@       @      3@              @       @     �N@      @      B@      @      @@       @      :@              @       @      @       @      9@      �?      @      �?      3@              @       @     �P@       @      M@      �?      =@      �?      ,@      �?      .@              =@              "@      �?      .@              Q@      3@      @@      0@      >@      $@      "@      $@      @      "@      @      �?      5@               @      @      B@      @      9@              &@      @      @       @      @      �?     �P@     @g@      N@     @g@      H@     �U@       @      <@      �?      9@      �?      @      G@      M@      .@      B@      .@      :@       @      :@      @      @      @      5@      �?      @      @      .@      @                      $@      ?@      6@      &@      0@      @       @       @       @      @       @      @      @      4@      @      (@      �?       @      @      @      @      @      �?      (@      Y@      �?      S@      �?      2@      �?      @              *@              M@      &@      8@      �?      3@      �?      @              ,@      $@      @      @      @      @       @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�>D5hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKkhth)h,K ��h.��R�(KKk��h{�B�         
                    @Dl���v�?�           @�@       @                           �?��<b���?             G@    r�                          ���3@�����H�?	             2@       ������������������������       �                     "@rm   rr������������������������       ��<ݚ�?             "@      D@       	                    @����X�?             <@     4@                          �4@�X�<ݺ?	             2@      0@������������������������       �r�q��?             @        ������������������������       �                     (@      $@������������������������       ��z�G��?             $@               N                    �?D��J<��?�           Є@      @       #                     �?���2���?!           �|@      �?                           �?uvI��?B            �X@      @                          �9@     ��?,             P@        ������������������������       �                     @      3@                           �?��Q:��?(            �M@     "@                           K@r�qG�?!             H@                                 �?��J�fj�?            �B@                                  ?@������?
             1@      ������������������������       ��C��2(�?             &@w      ������������������������       �      �?             @n                                �A@���Q��?             4@       ������������������������       �X�<ݚ�?             "@�      ������������������������       ����!pc�?             &@�                                �N@�C��2(�?             &@       ������������������������       �                     @c      ������������������������       �r�q��?             @      ������������������������       ��eP*L��?             &@             "                   @G@�ʻ����?             A@                                 �?����X�?             5@       ������������������������       ��<ݚ�?             "@V              !                   �@@�q�q�?
             (@       ������������������������       �      �?             @3      ������������������������       �      �?              @A      ������������������������       ��	j*D�?             *@�       $       -                    �?x�w�,�?�            pv@        %       &                   �7@��܂O�?1            �V@        ������������������������       �X�Cc�?	             ,@j       '       ,                   �=@�䞠�l�?(            @S@       (       +                    �?f>�cQ�?             �N@       )       *                 ���@�L���?            �B@        ������������������������       �                     &@�       ������������������������       �ȵHPS!�?             :@$       ������������������������       �      �?             8@       ������������������������       �                     0@       .       3                   �0@T�P*�/�?�            �p@        /       0                    $@8����?             7@        ������������������������       �և���X�?             @�       1       2                    �?      �?
             0@       ������������������������       �X�<ݚ�?             "@�       ������������������������       �                     @�       4       K                   �*@���0���?�            �n@       5       J                    �?4z�_�\�?|            �g@       6       ;                     @xP�Fֺ�?v            @f@       7       8                 `f�)@�����H�?            �F@        ������������������������       ��X�<ݺ?
             2@`      9       :                   �;@PN��T'�?             ;@       ������������������������       �                     ,@;      ������������������������       ��	j*D�?	             *@?      <       A                    7@��F���?\            �`@       =       >                 �?�@�?�|�?            �B@       ������������������������       �                     4@G       ?       @                   �3@�IєX�?             1@      ������������������������       ������H�?             "@!      ������������������������       �                      @�      B       I                 ���!@r�q��?D             X@      C       D                 ��@ ��~���?@            �V@        ������������������������       �և���X�?             @8      E       F                   �E@�gc� �?<            �T@      ������������������������       �ףp=
�?3            �Q@-      G       H                 P�@�θ�?	             *@      ������������������������       �                     @�      ������������������������       �      �?             @�       ������������������������       �      �?             @�       ������������������������       ��C��2(�?             &@v      L       M                 0��G@�h����?$             L@      ������������������������       �                     G@�      ������������������������       �ףp=
�?             $@�      O       X                     @��eN_:�?�             j@      P       U                    �? �^�@̩?J             ]@      Q       T                   �;@�����?>             W@        R       S                   �8@Pa�	�?            �@@      ������������������������       �                     9@-      ������������������������       �      �?              @%      ������������������������       �        )            �M@g      V       W                 ���`@�8��8��?             8@       ������������������������       �                     1@y       ������������������������       �����X�?             @}       Y       \                    �?��MΖ��??            @W@        Z       [                   �5@l��
I��?             ;@        ������������������������       �և���X�?             @        ������������������������       �      �?             4@        ]       d                    �?���|���?*            �P@       ^       _                    5@��
P��?            �A@        ������������������������       �                     @        `       c                    �?���Q��?             >@       a       b                   �@b�2�tk�?             2@        ������������������������       �      �?              @        ������������������������       ����Q��?             $@        ������������������������       ��q�q�?             (@        e       h                    �?�n`���?             ?@        f       g                    �?�q�q�?	             (@       ������������������������       ��q�q�?             @        ������������������������       �                     @        i       j                    @�KM�]�?
             3@       ������������������������       �                     &@        ������������������������       �      �?              @        �t�bh�h)h,K ��h.��R�(KKkKK��h\�B�        {@     `q@      $@      B@       @      0@              "@       @      @       @      4@      �?      1@      �?      @              (@      @      @     �z@     @n@     0w@     �U@     �N@     �B@      E@      6@      @             �B@      6@      ?@      1@      5@      0@      *@      @      $@      �?      @      @       @      (@      @      @      @       @      $@      �?      @              @      �?      @      @      3@      .@      .@      @      @       @       @      @      @      �?      @      @      @      "@     `s@     �H@     @R@      2@      @      "@      Q@      "@      J@      "@      A@      @      &@              7@      @      2@      @      0@             �m@      ?@      0@      @      @      @      (@      @      @      @      @             �k@      8@     �d@      7@     �c@      6@      D@      @      1@      �?      7@      @      ,@              "@      @      ]@      1@      B@      �?      4@              0@      �?       @      �?       @              T@      0@     @S@      *@      @      @     @R@      $@     �O@      @      $@      @      @              @      @      @      @      $@      �?     �K@      �?      G@              "@      �?     �J@     �c@      @     @\@      �?     �V@      �?      @@              9@      �?      @             �M@       @      6@              1@       @      @      I@     �E@       @      3@      @      @      @      .@      E@      8@      1@      2@      @              (@      2@      @      &@      �?      @      @      @      @      @      9@      @       @      @       @      @      @              1@       @      &@              @       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ���&hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKuhth)h,K ��h.��R�(KKu��h{�B@         V                    �?T�����?�           @�@      @       	                    $@R]�M2��?,           0}@ �<	�                             �?��a�n`�?             ?@ ��	�  ������������������������       �                     @�-}��                            �;@ �o_��?             9@      �?������������������������       �                     *@       @                           �?�q�q�?             (@      @������������������������       �����X�?             @      @������������������������       ����Q��?             @     �H@
       #                     �?Rԅ5l�?           @{@      "@                          �J@U��
�?=            @W@     @                        ��I/@և���X�?0            @S@      @������������������������       �                     @      8@                        ��";@r�q��?,             R@      �?������������������������       �z�G�z�?             $@      1@                           �?�U���?&             O@     �?                          �>@P����?             C@                                 �=@��S���?             .@       ������������������������       ��q�q�?             "@�      ������������������������       ��q�q�?             @w                              @��O@��<b���?             7@       ������������������������       �                      @�                                 �?�q�q�?
             .@       ������������������������       ��q�q�?             @�      ������������������������       ��q�q�?             "@�                                 �?      �?             8@       ������������������������       �                     @                                dT@�q�q�?             2@      ������������������������       ��eP*L��?             &@�      ������������������������       �؇���X�?             @(                                  M@      �?             0@       ������������������������       �                     @J      !       "                 `fF<@"pc�
�?	             &@       ������������������������       �                     @A      ������������������������       ��q�q�?             @�       $       S                 �T�I@��Z��?�            pu@       %       L                   �*@8d-���?�            �t@       &       +                 ���@��̋���?�            �n@        '       (                    �?�nkK�?             7@        ������������������������       �                      @�       )       *                   �:@��S�ۿ?             .@        ������������������������       �z�G�z�?             @�       ������������������������       �                     $@$       ,       -                   �1@,�(VB�?�            �k@        ������������������������       �և���X�?             @       .       ?                 ��L@@mW���?�            �j@        /       <                 ��@��ga�=�?.            �P@       0       3                   �8@PN��T'�?&             K@        1       2                 �Y�@�q�q�?
             (@        ������������������������       �z�G�z�?             @�       ������������������������       �                     @�       4       5                 ���@�����?             E@        ������������������������       �                     @�       6       7                 �Y�@(N:!���?            �A@       ������������������������       �"pc�
�?             &@�       8       9                  ��@�8��8��?             8@       ������������������������       �                     "@:      :       ;                   �<@�r����?
             .@      ������������������������       �                      @?      ������������������������       �����X�?             @I      =       >                 �?$@��
ц��?             *@       ������������������������       �����X�?             @G       ������������������������       ��q�q�?             @      @       G                 `f�)@�����?Z            `b@      A       B                     @�[|x��?K            �_@       ������������������������       �                     2@�      C       F                    �?h�WH��??             [@       D       E                 @!@ףp=
�?;             Y@      ������������������������       �l{��b��?0            �S@      ������������������������       ���s����?             5@-      ������������������������       �                      @,      H       I                   �;@��s����?             5@       ������������������������       �                      @�       J       K                   @B@�	j*D�?	             *@       ������������������������       �      �?              @v      ������������������������       �                     @�      M       N                    �?�d���?4            �U@       ������������������������       �                     1@�      O       P                    ?@��?^�k�?)            �Q@       ������������������������       �                     A@�      Q       R                   �A@�X�<ݺ?             B@        ������������������������       �����X�?             @      ������������������������       �                     =@-      T       U                    �?�q�q�?	             (@      ������������������������       �r�q��?             @g      ������������������������       �                     @�       W       `                     @^������?�            �n@       X       ]                 ���a@P���Q�?P             ^@       Y       \                    6@p� V�?G            �Y@        Z       [                   �/@@4և���?             <@       ������������������������       �                     3@        ������������������������       ��<ݚ�?             "@        ������������������������       �        5            �R@        ^       _                   �8@������?	             1@       ������������������������       �؇���X�?             @        ������������������������       ��z�G��?             $@        a       b                    @z�m�(�?D            @_@        ������������������������       ��q�q�?             (@        c       d                    -@3k���?<            @\@        ������������������������       �                     &@        e       p                    �?h+�v:�?7            �Y@       f       k                   �;@N1���?#            �N@       g       j                 ��@`՟�G��?             ?@        h       i                    �?������?	             .@       ������������������������       ����Q��?             $@        ������������������������       �                     @        ������������������������       �      �?	             0@        l       o                    �?d��0u��?             >@       m       n                 ���@      �?             2@        ������������������������       ����Q��?             @        ������������������������       ���
ц��?             *@        ������������������������       �r�q��?             (@        q       r                    �?���� �?            �D@        ������������������������       �և���X�?             @        s       t                 `fV6@������?             A@       ������������������������       ����Q��?             4@        ������������������������       �                     ,@        �t�bh�h)h,K ��h.��R�(KKuKK��h\�BP       0|@     Pp@     �v@      Y@      @      8@              @      @      2@              *@      @      @      @       @       @      @     �v@      S@      M@     �A@      F@     �@@      @             �C@     �@@       @       @     �B@      9@      9@      *@      @       @      @      @      @       @      2@      @       @              $@      @      @       @      @      @      (@      (@      @              @      (@      @      @      �?      @      ,@       @      @              "@       @      @              @       @     �r@     �D@     pr@      B@     @j@      A@      6@      �?       @              ,@      �?      @      �?      $@             �g@     �@@      @      @      g@      =@      J@      .@      G@       @       @      @      �?      @      @              C@      @      @              ?@      @      "@       @      6@       @      "@              *@       @       @              @       @      @      @       @      @      @       @     �`@      ,@      ]@      $@      2@             �X@      $@     �V@      $@     @R@      @      1@      @       @              1@      @       @              "@      @      @      @      @             @U@       @      1@              Q@       @      A@              A@       @      @       @      =@              @      @      �?      @      @              U@      d@      @     �\@       @     @Y@       @      :@              3@       @      @             �R@      @      *@      �?      @      @      @     �S@     �G@      @       @     �R@     �C@      &@             �O@     �C@     �@@      <@      ,@      1@      @      &@      @      @              @      $@      @      3@      &@      "@      "@       @      @      @      @      $@       @      >@      &@      @      @      :@       @      (@       @      ,@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�EhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKohth)h,K ��h.��R�(KKo��h{�B�         N                    �? ��ʀ_�?�           @�@      @                           @ʰ-M���?1           `~@ onal pr                        @3�4@�<ݚ�?             2@ o. 5: 2������������������������       �                     @ �.lib/p                           @���|���?	             &@       @������������������������       �                     @       @������������������������       �z�G�z�?             @      (@       ;                 ��i=@|������?#           @}@       	       :                 `f�:@��E�B��?�            �w@    �D@
                            �?���6�q�?�            �v@                                ��$:@������?             .@     �@@������������������������       �                     @       @������������������������       �      �?              @      @                            @0��QQX�?�            �u@       @                        `f�)@�Zl�i��?.            @T@       @������������������������       �                     @@      ,@                           �?ZՏ�m|�?             �H@       ������������������������       ����Q��?             @�                                �?@��2(&�?             F@       ������������������������       �                     1@w                                �*@�<ݚ�?             ;@       ������������������������       �      �?              @�                                 �?�KM�]�?
             3@      ������������������������       �                     &@�      ������������������������       �      �?              @�             3                   @@@(��R%��?�            �p@             0                   �<@BБ�|o�?}             j@                              ��@L(ݧa��?o             f@       ������������������������       �      �?             $@�             '                   �;@3��e��?i            �d@              &                   �3@4�{Y���?4            �T@              %                   �8@>A�F<�?0             S@      !       "                   �2@ �Cc}�?%             L@       ������������������������       �        
             ,@A      #       $                    �?؇���X�?             E@        ������������������������       ����Q��?             @�       ������������������������       ��L���?            �B@v       ������������������������       ����Q��?             4@j       ������������������������       �                     @�       (       +                 ��) @���N8�?5             U@       )       *                    �?p���?"             I@        ������������������������       ��C��2(�?             &@�       ������������������������       �                    �C@$       ,       -                    �?l��\��?             A@       ������������������������       ������H�?
             2@       .       /                    �?      �?	             0@       ������������������������       �ףp=
�?             $@]       ������������������������       �                     @�       1       2                   �?@     ��?             @@       ������������������������       �X�<ݚ�?             2@�       ������������������������       �d}h���?             ,@�       4       9                    �?���U�?(            �L@       5       6                   @C@`�q�0ܴ?!            �G@        ������������������������       �                     1@      7       8                 �?�@��S�ۿ?             >@       ������������������������       �                     1@`      ������������������������       �8�Z$���?
             *@:      ������������������������       �                     $@;      ������������������������       �        	             ,@?      <       K                    �?�x�(��?:             W@      =       B                    �?�ʻ����?.             Q@       >       A                   �@@\X��t�?             7@       ?       @                 0�&C@��S���?             .@       ������������������������       �և���X�?             @!      ������������������������       �      �?              @�      ������������������������       �      �?              @�      C       D                   �>@F�����?            �F@        ������������������������       ��<ݚ�?             "@8      E       J                     �?�E��ӭ�?             B@      F       G                    �?r�q��?             8@       ������������������������       �        	             &@,      H       I                    D@�	j*D�?	             *@      ������������������������       ��q�q�?             @�       ������������������������       �                     @�       ������������������������       �      �?             (@v      L       M                    @ �q�q�?             8@       ������������������������       �؇���X�?             @�      ������������������������       �                     1@�      O       l                    @f�z1�9�?�            @l@      P       U                    �?b��K�?�             j@       Q       T                    �?@4և���?             L@       R       S                 `�@1@������?            �B@       ������������������������       ����|���?             &@-      ������������������������       �                     :@%      ������������������������       �        
             3@g      V       k                    @J�V2���?k             c@       W       \                 `f�%@������?f             b@        X       Y                    �?
;&����?              G@        ������������������������       ��t����?             1@�       Z       [                 ��@J�8���?             =@        ������������������������       �����X�?             @        ������������������������       ��GN�z�?             6@        ]       b                    �?fhK�4�?F            �X@        ^       a                   �,@@�E�x�?!            �H@        _       `                   �;@�X�<ݺ?             2@        ������������������������       �      �?             @        ������������������������       �        	             ,@        ������������������������       �                     ?@        c       h                 039@`�Q��?%             I@        d       g                    �?ҳ�wY;�?             1@       e       f                 @3�/@�eP*L��?             &@        ������������������������       �      �?             @        ������������������������       �����X�?             @        ������������������������       �r�q��?             @        i       j                    �?6YE�t�?            �@@       ������������������������       �                     9@        ������������������������       �      �?              @        ������������������������       �      �?              @        m       n                    6@�t����?	             1@       ������������������������       �                      @        ������������������������       ��<ݚ�?             "@        �t�bh�h)h,K ��h.��R�(KKoKK��h\�B�       �|@     �o@     �x@     @W@      @      ,@              @      @      @              @      @      �?     Px@     �S@     �t@      H@     �s@      H@      &@      @      @              @      @     �r@      F@     @R@       @      @@             �D@       @      @       @      C@      @      1@              5@      @      @      @      1@       @      &@              @       @     �l@      B@     �e@      A@     @c@      7@      @      @     �b@      2@     @Q@      ,@      O@      ,@      I@      @      ,@              B@      @       @      @      A@      @      (@       @      @              T@      @     �H@      �?      $@      �?     �C@              ?@      @      0@       @      .@      �?      "@      �?      @              5@      &@      $@       @      &@      @     �K@       @     �F@       @      1@              <@       @      1@              &@       @      $@              ,@             �N@      ?@      C@      >@      $@      *@       @      @      @      @      @      @       @      @      <@      1@       @      @      :@      $@      4@      @      &@              "@      @       @      @      @              @      @      7@      �?      @      �?      1@             @P@      d@      I@     �c@      @      J@      @     �@@      @      @              :@              3@      G@     �Z@     �D@      Z@      8@      6@      @      (@      3@      $@       @      @      1@      @      1@     �T@      �?      H@      �?      1@      �?      @              ,@              ?@      0@      A@      &@      @      @      @      �?      @      @       @      @      �?      @      <@              9@      @      @      @      @      .@       @       @              @       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ4�phG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKahth)h,K ��h.��R�(KKa��h{�B@         &                     @@?�p�?�           @�@       @                           �?(�ruX��?�            0s@�                           �?rl[غ��?�            `k@��	�         	                 ��$:@�L�w��?U            �a@ l;�`f�l                           �?�IєX�?)             Q@                                 �J@���J��?"            �I@       ������������������������       �                    �G@      7@������������������������       �      �?             @      ,@������������������������       �@�0�!��?             1@      @
                         	>@ޚ)�?,             R@      @                        ��=@���>4��?             <@     @������������������������       �     ��?	             0@        ������������������������       ��q�q�?             (@       @                          �;@���!pc�?             F@                                  �7@      �?             $@      ?@������������������������       �                     @      @������������������������       �                     @Z                                 H@H�V�e��?             A@                                 �?H%u��?             9@       ������������������������       �                     $@w                              ��G@z�G�z�?             .@       ������������������������       ��q�q�?             @�      ������������������������       ������H�?             "@�      ������������������������       �X�<ݚ�?             "@�                              ��*@�Fǌ��?6            �S@                                 �9@�}�+r��?             3@       ������������������������       �z�G�z�?             @      ������������������������       �                     ,@      ������������������������       �        &             N@�             %                 `fmj@N�zv�?2             V@             $                    �?��Sݭg�?-            �S@               !                    2@�\��N��?             C@       ������������������������       �                     0@3      "       #                 03�R@�C��2(�?             6@      ������������������������       �        	             .@�       ������������������������       �����X�?             @�       ������������������������       �                     D@v       ������������������������       �      �?             $@j       '       L                    �?���iz�?�            Py@       (       G                 ��T?@P�I;l�?�            �q@       )       F                    �?țu���?�            @p@       *       C                    �?�*�w�?�             n@       +       >                   @@@�:�^���?�             l@       ,       /                    �?N�hƇ�?p             f@        -       .                   �7@ �o_��?             9@        ������������������������       �X�<ݚ�?             "@-       ������������������������       �      �?             0@]       0       3                 ���@�˹�m��?_             c@        1       2                    6@z�G�z�?	             .@        ������������������������       �                     @�       ������������������������       �      �?              @�       4       =                   �<@`�BX�l�?V             a@       5       <                 @3�@ ����?I            �]@       6       7                    �?(;L]n�?%             N@       ������������������������       �                     &@�       8       ;                   �5@@9G��?            �H@       9       :                 �?$@�����H�?             2@       ������������������������       �                     @;      ������������������������       �r�q��?             (@?      ������������������������       �                     ?@I      ������������������������       �        $            �M@7      ������������������������       �b�2�tk�?             2@G       ?       @                   �E@@��8��?             H@      ������������������������       �                     <@!      A       B                 P�@P���Q�?
             4@      ������������������������       �                     *@�      ������������������������       �؇���X�?             @8       D       E                    7@     ��?             0@      ������������������������       ��<ݚ�?             "@      ������������������������       �                     @-      ������������������������       �        
             3@,      H       I                    �?�û��|�?             7@       ������������������������       �X�<ݚ�?             "@�       J       K                 ���E@����X�?	             ,@        ������������������������       �և���X�?             @v      ������������������������       �                     @�      M       Z                    �?Υf���?D            �^@      N       S                    7@Z��Yo��?$             O@       O       P                    0@l��[B��?             =@       ������������������������       �r�q��?             (@�      Q       R                 ��!@������?             1@        ������������������������       �      �?             @      ������������������������       ��C��2(�?             &@-      T       Y                    �?r٣����?            �@@      U       X                    =@����X�?             5@      V       W                  ��@r�q��?
             (@       ������������������������       �                      @y       ������������������������       �      �?             @}       ������������������������       �X�<ݚ�?             "@�       ������������������������       �r�q��?             (@        [       `                 03�9@�0u��A�?              N@       \       _                    @d�
��?             F@       ]       ^                    �?��.k���?             A@        ������������������������       �r�q��?             (@        ������������������������       ����|���?             6@        ������������������������       �      �?             $@        ������������������������       �        
             0@        �t�bh�h)h,K ��h.��R�(KKaKK��h\�B       �{@     �p@      a@     @e@      \@     �Z@     �[@      =@      P@      @      I@      �?     �G@              @      �?      ,@      @     �G@      9@      .@      *@      &@      @      @       @      @@      (@      @      @      @                      @      ;@      @      6@      @      $@              (@      @      @       @       @      �?      @      @      �?     �S@      �?      2@      �?      @              ,@              N@      9@     �O@      4@      M@      4@      2@              0@      4@       @      .@              @       @              D@      @      @     0s@     �X@     �n@      B@      m@      ;@     �j@      ;@     �i@      4@     �c@      3@      2@      @      @      @      ,@       @     �a@      (@      (@      @      @              @      @      `@      "@     @]@       @      M@       @      &@             �G@       @      0@       @      @              $@       @      ?@             �M@              &@      @     �G@      �?      <@              3@      �?      *@              @      �?      "@      @       @      @      @              3@              ,@      "@      @      @      $@      @      @      @      @              N@      O@      7@     �C@      .@      ,@       @      $@      *@      @      @      @      $@      �?       @      9@      @      .@       @      $@               @       @       @      @      @       @      $@     �B@      7@      5@      7@      0@      2@       @      $@      ,@       @      @      @      0@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJLxhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK
hsKahth)h,K ��h.��R�(KKa��h{�B@         N                 0�^I@^IB�A��?�           @�@      @                         �#@�q�q��?n            �@ �ژ�                          ���@�����=�?�            0p@�y��                             �?V�L��?X            �`@#y��                          ��@ ˤ���?H            �Z@              	                   �:@xdQ�m��?7            @T@      @                        ��@��2(&�?             6@      ,@������������������������       ����!pc�?             &@      2@������������������������       �        	             &@       @
                           �?���#�İ?&            �M@      B@                          �=@HP�s��?             9@     3@������������������������       ������H�?             2@      (@������������������������       �                     @      "@������������������������       �                     A@       @������������������������       �$��m��?             :@        ������������������������       ��<ݚ�?             ;@                                  �:@�ص�ݒ�?N            @_@                                  �?`2U0*��?             I@      ������������������������       �                    �B@�      ������������������������       �8�Z$���?             *@w                                 �?��n�?1            �R@       ������������������������       ����Q��?             @�                              �?�@b�h�d.�?-            �Q@       ������������������������       �        
             ,@�                                @@@d}h���?#             L@      ������������������������       �r֛w���?             ?@c                              pf� @�J�4�?             9@      ������������������������       �z�G�z�?             .@      ������������������������       �ףp=
�?             $@�             5                    �?��2X�K�?�            �s@             $                    �?@S�)�q�?t            �f@               !                     �?�q�q�?             5@       ������������������������       �                     @3      "       #                    ;@��S���?
             .@       ������������������������       �      �?             @�       ������������������������       ����|���?             &@�       %       0                    �?�Zű���?e             d@       &       /                    �?X�;�^o�?F            �[@       '       *                     �?�T|n�q�?8            �U@        (       )                 `f�;@      �?             <@       ������������������������       �p�ݯ��?             3@�       ������������������������       �                     "@�       +       .                     @�y��*�?&             M@       ,       -                    5@���c���?"             J@        ������������������������       �����X�?             @       ������������������������       ������H�?            �F@-       ������������������������       �                     @]       ������������������������       �                     8@�       1       4                    $@d,���O�?            �I@        2       3                    @�E��ӭ�?             2@       ������������������������       �                     (@�       ������������������������       �r�q��?             @�       ������������������������       �                    �@@�       6       K                    @� Mv:�?T            �`@      7       J                    @HC>���?L            �^@       8       A                     @L���a��?F            �\@      9       @                    �?����e��?)            �P@      :       ;                     �?��Y��]�?            �D@       ������������������������       �                     @?      <       ?                   �*@г�wY;�?             A@      =       >                 ��Y)@�X�<ݺ?             2@       ������������������������       �                     "@G       ������������������������       ������H�?             "@      ������������������������       �                     0@!      ������������������������       �                     9@�      B       E                    �?f�Sc��?            �H@       C       D                  S�-@��s����?             5@        ������������������������       �z�G�z�?             @8      ������������������������       �        	             0@      F       I                    :@      �?             <@      G       H                    ,@�n_Y�K�?	             *@       ������������������������       �      �?             @�      ������������������������       ��q�q�?             "@�       ������������������������       ����Q��?             .@�       ������������������������       �և���X�?             @v      L       M                    !@8�Z$���?             *@       ������������������������       ��q�q�?             @�      ������������������������       �                     @�      O       Z                   �=@�g+�v�?V             a@       P       Y                    @�5��?%             K@      Q       V                    �?���Q �?             �H@        R       U                   �;@
j*D>�?             :@      S       T                   �8@ҳ�wY;�?             1@      ������������������������       ����Q��?             $@%      ������������������������       �                     @g      ������������������������       �                     "@�       W       X                 83G`@���}<S�?             7@       ������������������������       �        	             ,@}       ������������������������       ��<ݚ�?             "@�       ������������������������       �                     @        [       `                    �?R�(CW�?1            �T@        \       _                    �?h+�v:�?             A@        ]       ^                  �	U@����X�?             ,@        ������������������������       �      �?              @        ������������������������       �r�q��?             @        ������������������������       ��G�z��?             4@        ������������������������       �                     H@        �t�bh�h)h,K ��h.��R�(KKaKK��h\�B       �z@     �q@     `x@     @g@      j@     �I@     �X@     �A@     @W@      ,@      S@      @      3@      @       @      @      &@             �L@       @      7@       @      0@       @      @              A@              1@      "@      @      5@     @[@      0@      H@       @     �B@              &@       @     �N@      ,@      @       @      M@      (@      ,@              F@      (@      7@       @      5@      @      (@      @      "@      �?     �f@     �`@     �b@      A@      ,@      @      @               @      @      �?      @      @      @     �`@      ;@      X@      ,@      R@      ,@      5@      @      (@      @      "@             �I@      @     �F@      @      @       @      D@      @      @              8@              C@      *@      @      *@              (@      @      �?     �@@              A@     @Y@      7@     �X@      3@      X@      �?     @P@      �?      D@              @      �?     �@@      �?      1@              "@      �?       @              0@              9@      2@      ?@      @      1@      @      �?              0@      ,@      ,@      @       @       @       @      @      @      "@      @      @      @      &@       @      @       @      @             �A@     @Y@      6@      @@      1@      @@      .@      &@      @      &@      @      @              @      "@               @      5@              ,@       @      @      @              *@     @Q@      *@      5@      @      $@      @      @      �?      @      "@      &@              H@�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJW��8hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKshth)h,K ��h.��R�(KKs��h{�B�         L                    �?��!h
��?�           @�@      @                           @>���_�?           �{@ �B	�                             @�q�q�?             2@0��  ������������������������       �                     &@�����  ������������������������       �؇���X�?             @       @                            �?$���'w�?           �z@                                  @C@���%&�?3            �S@     @                           �?      �?             E@     @	                          �?@)O���?             B@     @
                        `f�N@��}*_��?             ;@     @������������������������       �և���X�?             5@      @������������������������       �r�q��?             @        ������������������������       ��<ݚ�?             "@      �?������������������������       ��q�q�?             @      X@                           @@���"͏�?            �B@     �@@                          �F@�q�q�?
             (@      0@������������������������       �      �?             @Z      ������������������������       ��q�q�?             @�                                 �?�J�4�?             9@       ������������������������       �                     $@w                              03�S@������?	             .@       ������������������������       �      �?              @�      ������������������������       �                     @�             ?                    @@������?�            �u@             >                    @��ē*�?�            pp@                                 �?��]��?�            @o@                               �2@���?            �D@                                @@:ɨ��?            �@@      ������������������������       ��S����?             3@�      ������������������������       �      �?             ,@(      ������������������������       �                      @V              ;                    �?� ����?�             j@      !       :                   �?@L(ݧa��?n             f@      "       7                   �<@|T(W�j�?g            �d@      #       (                     @�8��8��?\             b@        $       %                    @�����H�?             B@        ������������������������       �                     @v       &       '                    5@�r����?             >@        ������������������������       �z�G�z�?             $@�       ������������������������       �ףp=
�?             4@�       )       *                 ��@�>����?F             [@        ������������������������       �      �?              @�       +       6                 pf� @ "��u�?A             Y@       ,       3                 @3�@�˹�m��?3             S@       -       .                    �?�nkK�?#             G@        ������������������������       �؇���X�?             @-       /       2                 ��L@ ���J��?            �C@       0       1                    :@P���Q�?             4@       ������������������������       �        	             *@A       ������������������������       �؇���X�?             @�       ������������������������       �                     3@�       4       5                   �4@�r����?             >@        ������������������������       ����|���?             &@�       ������������������������       �                     3@      ������������������������       �                     8@�       8       9                   �=@��s����?             5@       ������������������������       �      �?              @:      ������������������������       �$�q-�?             *@;      ������������������������       ��q�q�?             (@?      <       =                    6@     ��?             @@      ������������������������       ������?             5@7      ������������������������       ����|���?             &@G       ������������������������       �        	             *@      @       K                   �M@ 	��p�?8            �U@      A       J                   �*@xdQ�m��?4            @T@      B       I                   `F@0��_��?"            �J@      C       H                 `fF)@�ݜ�?            �C@       D       E                 �?�@��S�ۿ?             >@       ������������������������       �        	             ,@      F       G                    C@      �?             0@      ������������������������       �                      @,      ������������������������       �      �?              @�      ������������������������       ��q�q�?             "@�       ������������������������       �        	             ,@�       ������������������������       �                     <@v      ������������������������       �r�q��?             @�      M       r                    @Ȩ�I��?�            �p@      N       Y                     @��yn�?�            p@      O       T                   �;@ 7���B�?Q            �`@       P       Q                   �7@���}<S�?             G@      ������������������������       �                    �@@�       R       S                    �?�	j*D�?             *@       ������������������������       �      �?              @-      ������������������������       ����Q��?             @%      U       X                 03�>@ }�Я��?6            @V@       V       W                   �H@P�Lt�<�?             C@       ������������������������       �                     <@y       ������������������������       �ףp=
�?             $@}       ������������������������       �                    �I@�       Z       g                   �9@��\j���?H            �^@        [       \                  s�@>4և���?!             L@        ������������������������       �                     @        ]       b                    �?�J��%�?            �H@       ^       a                    �?П[;U��?             =@       _       `                 �&B@��H�}�?             9@        ������������������������       ����Q��?             @        ������������������������       ��z�G��?             4@        ������������������������       �                     @        c       d                    @R���Q�?             4@        ������������������������       �      �?             @        e       f                    3@      �?	             0@       ������������������������       �                     $@        ������������������������       �r�q��?             @        h       q                 ��Y7@���|���?'            �P@       i       p                   @B@�c�Α�?#             M@       j       m                    �?z�G�z�?             I@       k       l                   �;@r٣����?            �@@        ������������������������       �                     "@        ������������������������       ��q�q�?             8@        n       o                   �0@�t����?	             1@       ������������������������       �      �?              @        ������������������������       �                     "@        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                      @        �t�b�       h�h)h,K ��h.��R�(KKsKK��h\�B0       �z@     �q@     �v@     �U@      @      (@              &@      @      �?      v@     �R@     �H@      >@      5@      5@      3@      1@      1@      $@      (@      "@      @      �?       @      @       @      @      <@      "@      @      @      @      @      @       @      5@      @      $@              &@      @      @      @      @             s@     �F@      l@     �C@     `j@     �C@      ?@      $@      7@      $@      0@      @      @      @       @             �f@      =@     @c@      7@     �b@      0@     �`@      (@      @@      @      @              :@      @       @       @      2@       @      Y@       @      @       @     �W@      @     �Q@      @      F@       @      @      �?      C@      �?      3@      �?      *@              @      �?      3@              :@      @      @      @      3@              8@              1@      @      @      @      (@      �?      @      @      :@      @      3@       @      @      @      *@             @T@      @      S@      @      H@      @      A@      @      <@       @      ,@              ,@       @       @              @       @      @      @      ,@              <@              @      �?     �Q@     `h@      O@     `h@      @     @`@      @      E@             �@@      @      "@       @      @       @      @      �?      V@      �?     �B@              <@      �?      "@             �I@     �L@     @P@     �@@      7@              @     �@@      0@      0@      *@      0@      "@       @      @      ,@      @              @      1@      @       @       @      .@      �?      $@              @      �?      8@      E@      0@      E@      $@      D@       @      9@              "@       @      0@       @      .@       @      @              "@      @       @       @               @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��UhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKhth)h,K ��h.��R�(KK��h{�B�         Z                    �?����?�           @�@     &@                           @���Ee�?6           p~@      .@                        @3�4@8����?             7@        ������������������������       �                     $@      @                            @��
ц��?
             *@        ������������������������       �                     @     �F@������������������������       �                     @      $@       U                 03�U@��2�
�?&            }@     =@	       <                 039@8�ƨxt�?           �{@     @
                           �?������?�            �t@       @                            @��k=.��?            �G@      @������������������������       �r�q��?             @      �?������������������������       �� ��1�?            �D@      @       +                   �<@h��=�?�            �q@     @       "                   �;@t��ճC�?p             f@     @                          �7@`�H�/��?D            �Y@     @                           �?@4և���?,            �Q@                                �3@�.ߴ#�?%            �N@                                  @�˹�m��?             C@       ������������������������       ������H�?             "@w                                �0@ 	��p�?             =@       ������������������������       �      �?              @�                              ��Y @���N8�?             5@      ������������������������       �ףp=
�?             $@�      ������������������������       �                     &@�      ������������������������       �                     7@c      ������������������������       ��<ݚ�?             "@                              �&B@     ��?             @@       ������������������������       �X�<ݚ�?             "@�             !                 ��)"@�nkK�?             7@                               �?�@�C��2(�?	             &@       ������������������������       �                     @J      ������������������������       �z�G�z�?             @3      ������������������������       �                     (@A      #       *                    �?�?�|�?,            �R@       $       %                     @��v$���?$            �N@        ������������������������       �                     $@v       &       '                    �?���J��?            �I@        ������������������������       �                     1@�       (       )                 ��) @г�wY;�?             A@       ������������������������       �                     9@�       ������������������������       ������H�?             "@�       ������������������������       �$�q-�?             *@$       ,       ;                    �?T>D5j�?E            @Z@       -       8                   @F@�+�$f��?@            �X@       .       7                 ��+@d1<+�C�?.            @R@       /       6                    D@     ��?(             P@       0       5                 `fF)@\-��p�?$             M@       1       2                   @@@ףp=
�?              I@        ������������������������       �z�G�z�?             4@�       3       4                   @C@(;L]n�?             >@       ������������������������       �                     9@�       ������������������������       �z�G�z�?             @�       ������������������������       �      �?              @      ������������������������       ��q�q�?             @�       ������������������������       �                     "@`      9       :                    M@`2U0*��?             9@      ������������������������       �                     4@;      ������������������������       �z�G�z�?             @?      ������������������������       �                     @I      =       D                 ��";@F�t�K��?F            �\@       >       A                 ��$:@���Q��?             9@        ?       @                   �@@�	j*D�?             *@       ������������������������       �      �?              @!      ������������������������       �                     @�      B       C                   �F@      �?             (@       ������������������������       �����X�?             @8       ������������������������       �z�G�z�?             @8      E       R                 03�M@4�<����?6            @V@      F       Q                    �?L=�m��?(            �N@      G       H                    �?��Hg���?            �F@       ������������������������       ��C��2(�?             &@�      I       P                    �?�t����?             A@       J       K                   @>@>���Rp�?             =@        ������������������������       ����Q��?             @v      L       O                 03�I@r�q��?             8@      M       N                 �T�@@�}�+r��?             3@       ������������������������       �؇���X�?             @�      ������������������������       �                     (@�      ������������������������       ����Q��?             @�      ������������������������       ����Q��?             @�       ������������������������       �        	             0@      S       T                    �?h�����?             <@      ������������������������       �P���Q�?	             4@%      ������������������������       �                      @g      V       Y                   �D@8�A�0��?             6@       W       X                    �?և���X�?	             ,@        ������������������������       ��q�q�?             @}       ������������������������       �      �?              @�       ������������������������       �      �?              @        [       ~                    @��PN���?�             l@       \       e                     @�E+]9��?�            `k@       ]       ^                    @��sK�z�?P            �^@        ������������������������       �և���X�?             @        _       d                 03[=@XB���?K             ]@        `       c                    :@�:�^���?            �F@       a       b                   �;@г�wY;�?             A@        ������������������������       ������H�?             "@        ������������������������       �                     9@        ������������������������       ����!pc�?             &@        ������������������������       �        /            �Q@        f       k                 �̌@r�q��?@             X@        g       j                    �?      �?             8@       h       i                 ���@r�q��?
             2@        ������������������������       �                      @        ������������������������       ��z�G��?             $@        ������������������������       �                     @        l       }                   @B@X�<ݚ�?1             R@       m       n                    @�g�y��?+             O@        ������������������������       �r�q��?             @        o       |                    �?~h����?&             L@       p       w                    �?z�):���?!             I@       q       t                    �?և���X�?             <@       r       s                   �;@j���� �?             1@       ������������������������       �      �?              @        ������������������������       ��<ݚ�?             "@        u       v                 @3�/@�eP*L��?             &@        ������������������������       �      �?             @        ������������������������       ����Q��?             @        x       y                   �9@�X����?             6@        ������������������������       �և���X�?             @        z       {                    �?������?	             .@        ������������������������       ������H�?             "@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KKKK��h\�B�        }@      o@     �y@     �S@      @      0@              $@      @      @              @      @             y@     �O@     @x@      K@     �r@      @@      C@      "@      @      �?     �@@       @      p@      7@     �d@      (@      W@      $@     @P@      @      M@      @     �A@      @       @      �?      ;@       @      @      �?      4@      �?      "@      �?      &@              7@              @       @      ;@      @      @      @      6@      �?      $@      �?      @              @      �?      (@              R@       @      N@      �?      $@              I@      �?      1@             �@@      �?      9@               @      �?      (@      �?     �W@      &@     �U@      &@     �O@      $@      K@      $@      I@       @     �F@      @      0@      @      =@      �?      9@              @      �?      @      @      @       @      "@              8@      �?      4@              @      �?      @              W@      6@      .@      $@      "@      @      @      @      @              @      @       @      @      @      �?     @S@      (@      I@      &@      A@      &@      $@      �?      8@      $@      6@      @       @      @      4@      @      2@      �?      @      �?      (@               @      @       @      @      0@              ;@      �?      3@      �?       @              *@      "@      @       @       @      @      @      @      @      �?      L@      e@      I@      e@      @      ]@      @      @      @      \@      @     �D@      �?     �@@      �?       @              9@      @       @             �Q@     �E@     �J@      @      5@      @      .@               @      @      @              @      D@      @@      >@      @@      �?      @      =@      ;@      7@      ;@      0@      (@      $@      @      @      @      @       @      @      @      @      @      @       @      @      .@      @      @      @      &@      �?       @      @      @      @              $@              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��DphG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK
hsK]hth)h,K ��h.��R�(KK]��h{�B@         4                    �?���x�W�?�           @�@     &@       	                 �?�@�.��q�?!           �|@ , 4.],                           @@@�\�)G�?Z            �`@ be use                           �?=�Ѝ;�?H            �Y@> x1 =                           �<@L�[2[
�?A            �V@     �?������������������������       �p`q�q��?;            �S@      �?������������������������       �      �?             (@      @������������������������       �      �?             (@        ������������������������       �                     @@      �?
       /                    �?�A����?�            �t@     �?                            �?��0�ϥ�?�            �q@      &@                           �?��H���?8            @Y@      @                          �>@*;L]n�?3            �V@                                   ?@<=�,S��?            �A@       ������������������������       ��G��l��?
             5@                                  �E@؇���X�?             ,@      @������������������������       ������H�?             "@Z      ������������������������       �z�G�z�?             @�                                 �?�2�o�U�?!            �K@                                  �?�g�y��?             ?@                              `��f@b�2�tk�?	             2@      ������������������������       ����!pc�?             &@�      ������������������������       �և���X�?             @�      ������������������������       ��	j*D�?             *@�                              ��yC@ �q�q�?             8@       ������������������������       �z�G�z�?             @c      ������������������������       �                     3@      ������������������������       ����|���?             &@                                  �?�0��D/�?w            �f@                                  �?��.k���?             1@      ������������������������       ��eP*L��?             &@V      ������������������������       ��q�q�?             @J      !       "                 @3�@�N˹|�?l            �d@       ������������������������       ��q�q�?             (@A      #       (                 м[3@n�3���?g             c@       $       '                    �?��.���?J            @\@       %       &                    �?�	��)��?C            �Y@       ������������������������       ��S����?=            �W@j       ������������������������       �                      @�       ������������������������       �z�G�z�?             $@�       )       ,                    �?��-�=��?            �C@        *       +                    ;@�}�+r��?             3@        ������������������������       �z�G�z�?             @$       ������������������������       �        
             ,@       -       .                     @R���Q�?             4@       ������������������������       ��z�G��?	             $@-       ������������������������       �                     $@]       0       3                   �C@���.�6�?             G@        1       2                 мK;@r�q��?             2@        ������������������������       �                     "@�       ������������������������       ��q�q�?             "@�       ������������������������       �                     <@�       5       >                     @
��l۹�?�             o@        6       7                    �?�8���?M             ]@       ������������������������       �                     9@�       8       =                   �;@���L��?<            �V@       9       :                    6@�n`���?             ?@       ������������������������       �      �?              @;      ;       <                    �?���}<S�?             7@      ������������������������       �                     .@I      ������������������������       �      �?              @7      ������������������������       �        %             N@G       ?       \                    B@B��仱�?V            �`@      @       U                    �?����v��?O            �^@      A       H                    �?�W*��?<            @X@       B       G                    �?p9W��S�?             C@      C       D                    �?     ��?             @@        ������������������������       �և���X�?             @8      E       F                 ��@ �o_��?             9@       ������������������������       ����Q��?             @-      ������������������������       �z�G�z�?
             4@,      ������������������������       �r�q��?             @�      I       T                    �?Ɣ��Hr�?$            �M@       J       Q                 `f�%@z�J��?            �G@       K       L                   �@R�}e�.�?             :@       ������������������������       �����X�?             @�      M       P                    �?�KM�]�?             3@      N       O                   �9@r�q��?	             (@       ������������������������       �                     @�      ������������������������       �����X�?             @�      ������������������������       �                     @�       R       S                    =@���N8�?             5@      ������������������������       ��r����?             .@-      ������������������������       �      �?             @%      ������������������������       �                     (@g      V       Y                    �?$��m��?             :@        W       X                   �9@�q�q�?             "@        ������������������������       �      �?             @}       ������������������������       ����Q��?             @�       Z       [                 ��p@@@�0�!��?             1@        ������������������������       �      �?              @        ������������������������       �                     "@        ������������������������       �ףp=
�?             $@        �t�bh�h)h,K ��h.��R�(KK]KK��h\�B�       P{@     0q@     `v@     @Z@     �^@      *@     �V@      *@     @T@      $@      R@      @      "@      @      "@      @      @@             �m@      W@      h@     @V@     �K@      G@     �I@     �C@      *@      6@      &@      $@       @      (@      �?       @      �?      @      C@      1@      .@      0@      &@      @       @      @      @      @      @      "@      7@      �?      @      �?      3@              @      @     @a@     �E@      "@       @      @      @      @       @      `@     �A@      @       @     @_@      ;@     �V@      7@      V@      .@      T@      .@       @               @       @     �A@      @      2@      �?      @      �?      ,@              1@      @      @      @      $@             �E@      @      .@      @      "@              @      @      <@             �S@     @e@      @     �[@              9@      @     @U@      @      9@      @      @       @      5@              .@       @      @              N@     @R@      N@      P@     �M@     �G@      I@      &@      ;@      $@      6@      @      @      @      2@      @       @      @      0@      �?      @      B@      7@      8@      7@      3@      @       @      @      1@       @      $@       @      @              @       @      @              @      0@       @      *@      @      @      (@              1@      "@      @      @      �?      @       @      @      ,@      @      @      @      "@              "@      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ%�[6hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKmhth)h,K ��h.��R�(KKm��h{�B@         T                    �?�25����?�           @�@     &@                           �?�NG�#=�?/           �}@     �;@                           +@�(~�[�?4            �U@      �?������������������������       �      �?              @      @                           �?�2��?0            �S@     0@                        ���@P̏����?             �L@      "@������������������������       �                     &@      @                        `f�B@8����?             G@      @	       
                 0C�;@*O���?             B@     7@������������������������       �8^s]e�?             =@       @������������������������       �և���X�?             @        ������������������������       �ףp=
�?             $@      @                          �9@�eP*L��?             6@        ������������������������       ����|���?             &@     @U@                           D@���!pc�?
             &@     .@������������������������       �                     @     �M@������������������������       �      �?             @                                   @n�i8�?�            px@                                   �?�X����?             6@                                   @������?
             .@        ������������������������       �                      @        ������������������������       �և���X�?             @        ������������������������       �և���X�?             @               #                     �?s�As��?�            w@                                   �>@�iޤ��?)            �P@                                 @D@�'�=z��?            �@@                                �̌/@������?
             .@        ������������������������       �                     @        ������������������������       ����Q��?             $@                                   K@�q�q�?             2@       ������������������������       �8�Z$���?             *@        ������������������������       �z�G�z�?             @        !       "                    �?�t����?             A@       ������������������������       �        	             ,@A      ������������������������       �z�G�z�?             4@�       $       Q                    �?|b�!]	�?�            �r@       %       ,                  ��@t�6Z���?�            0q@        &       '                 ��@���7�?             F@        ������������������������       �        
             2@�       (       )                    7@$�q-�?             :@        ������������������������       �                     (@�       *       +                 ���@؇���X�?
             ,@        ������������������������       ��q�q�?             @$       ������������������������       �                      @       -       4                   �:@4�^���?�            �l@        .       3                 ��Y @@�j;��?1            �Q@       /       0                   �4@b�h�d.�?            �A@        ������������������������       ��	j*D�?
             *@�       1       2                 P�N@�C��2(�?             6@        ������������������������       ����Q��?             @�       ������������������������       �                     1@�       ������������������������       �                     B@�       5       D                   @@@z�G�z�?h             d@       6       C                 039@�DC��,�?=            �V@      7       :                 pb@l������?6            �S@        8       9                 ��@b�2�tk�?             2@      ������������������������       ����!pc�?             &@:      ������������������������       �և���X�?             @;      ;       B                   �>@��.��?+            �N@      <       =                 pf� @$�q-�?%             J@       ������������������������       �                     9@7      >       ?                     @PN��T'�?             ;@        ������������������������       �      �?              @      @       A                    �?�KM�]�?             3@      ������������������������       �ףp=
�?             $@�      ������������������������       ������H�?             "@�      ������������������������       ��q�q�?             "@8       ������������������������       �      �?             (@8      E       P                   �J@�LQ�1	�?+            @Q@      F       O                   �F@X��Oԣ�?&             O@      G       H                 @3�@��0{9�?            �G@       ������������������������       �      �?             0@�      I       N                    �?��a�n`�?             ?@       J       M                     @H%u��?             9@       K       L                   @A@���!pc�?	             &@       ������������������������       ��q�q�?             @�      ������������������������       �z�G�z�?             @�      ������������������������       �                     ,@�      ������������������������       �                     @�      ������������������������       �        	             .@�      ������������������������       �����X�?             @�       R       S                    $@ 7���B�?             ;@       ������������������������       ������H�?             "@-      ������������������������       �                     2@%      U       ^                 `f�$@�<ݚ�?�            @m@       V       Y                    �?և���X�?%             L@        W       X                 ���@r�q��?             8@        ������������������������       �����X�?             @}       ������������������������       ��t����?             1@�       Z       ]                    ;@      �?             @@       [       \                 ���@r�q��?             8@        ������������������������       �                     @        ������������������������       �������?             1@        ������������������������       �      �?              @        _       d                     @4\�����?q            @f@       `       c                   �;@`���i��?P            �`@        a       b                   �8@t��ճC�?             F@       ������������������������       �                     C@        ������������������������       �      �?             @        ������������������������       �        3             V@        e       l                 `v�6@(옄��?!             G@       f       g                    @     ��?             @@        ������������������������       �                     @        h       i                 `�/@� �	��?             9@        ������������������������       �؇���X�?             @        j       k                    >@�E��ӭ�?             2@       ������������������������       ����|���?             &@        ������������������������       �؇���X�?             @        ������������������������       �        	             ,@        �t�bh�h)h,K ��h.��R�(KKmKK��h\�B�       pz@     r@     0w@     �Z@      L@      ?@      �?      @     �K@      8@     �E@      ,@      &@              @@      ,@      7@      *@      4@      "@      @      @      "@      �?      (@      $@      @      @       @      @      @              �?      @     �s@      S@      @      .@      @      &@               @      @      @      @      @     @s@     �N@     �G@      4@      1@      0@      &@      @      @              @      @      @      (@       @      &@      @      �?      >@      @      ,@              0@      @     Pp@     �D@     `m@      D@      E@       @      2@              8@       @      (@              (@       @      @       @       @              h@      C@     @P@      @      =@      @      "@      @      4@       @      @       @      1@              B@              `@      @@      Q@      7@      O@      1@      &@      @       @      @      @      @     �I@      $@      H@      @      9@              7@      @      @       @      1@       @      "@      �?       @      �?      @      @      @      @      N@      "@     �K@      @      D@      @      (@      @      <@      @      6@      @       @      @      @       @      @      �?      ,@              @              .@              @       @      :@      �?       @      �?      2@              J@     �f@      8@      @@      @      4@       @      @       @      .@      4@      (@      *@      &@              @      *@      @      @      �?      <@     �b@      @      `@      @     �D@              C@      @      @              V@      9@      5@      &@      5@              @      &@      ,@      @      �?      @      *@      @      @      �?      @      ,@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�	3 hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKqhth)h,K ��h.��R�(KKq��h{�B@         .                 `f�%@T�����?�           @�@      @                        ���@.�*���?�            �r@     �B@                        03s@�Ń��̧?             E@     @������������������������       �                     ?@      �?������������������������       ��C��2(�?             &@      &@       	                    �?ά��.��?�            @p@     �N@                        ���@�	j*D�?             :@        ������������������������       �X�<ݚ�?             "@      �?������������������������       �@�0�!��?             1@     �D@
       #                    �?P�G��l�?�            @m@      @                          �>@N���X�?n            �e@                                  �? d��u�?M            @_@     @                          �5@���^���?G            �\@                                   1@д>��C�?             =@      @������������������������       ��<ݚ�?             "@      @                        ��L@R���Q�?             4@       @������������������������       �      �?              @Z      ������������������������       ��8��8��?	             (@�                                �<@��+��<�?6            �U@                              P��@�(\����?2             T@       ������������������������       �      �?              @n                                �;@�k~X��?.             R@                                 �9@���N8�?             5@      ������������������������       �                     ,@�      ������������������������       �؇���X�?             @�      ������������������������       �                    �I@c      ������������������������       �r�q��?             @      ������������������������       ����Q��?             $@                              �&B@      �?!             H@       ������������������������       �        	             &@(                                 @@@4�B��?            �B@       ������������������������       �z�G�z�?             $@J      !       "                   �E@PN��T'�?             ;@      ������������������������       �                     .@A      ������������������������       ��q�q�?             (@�       $       %                 ���@�p����?%            �N@        ������������������������       �                     @v       &       '                    �?N{�T6�?!            �K@        ������������������������       ��q�q�?	             (@�       (       )                     @��V#�?            �E@        ������������������������       �                     @�       *       +                   �9@��Sݭg�?            �C@        ������������������������       ��t����?
             1@$       ,       -                    A@���|���?
             6@       ������������������������       ���
ц��?             *@       ������������������������       ��<ݚ�?             "@-       /       R                    �?\����?�            �y@       0       O                 Ј�V@�D�>��?�            �l@       1       N                    �?�϶O'3�?�            @j@       2       3                    ,@� $jS`�?r            �f@        ������������������������       �        
             *@�       4       ;                    �?B��Z��?h            @e@        5       6                  A7@*O���?             B@        ������������������������       �z�G�z�?             $@      7       :                   @B@���B���?             :@       8       9                    �?R���Q�?             4@      ������������������������       �z�G�z�?             .@:      ������������������������       �                     @;      ������������������������       ��q�q�?             @?      <       M                    �?��v����?S            �`@      =       D                 `fF:@�MI8d�?E            �[@      >       ?                    ?@0z�(>��?,            �Q@       ������������������������       �                    �F@      @       A                   �*@ȵHPS!�?             :@       ������������������������       �"pc�
�?             &@�      B       C                    �?��S�ۿ?             .@      ������������������������       �                     $@8       ������������������������       �z�G�z�?             @8      E       H                   �>@      �?             D@       F       G                   �J@����X�?             ,@       ������������������������       �r�q��?             @,      ������������������������       �      �?              @�      I       L                     @���B���?             :@       J       K                    @@�}�+r��?             3@       ������������������������       ������H�?             "@v      ������������������������       �                     $@�      ������������������������       �և���X�?             @�      ������������������������       �                     7@�      ������������������������       �                     ;@�      P       Q                    �?�\��N��?
             3@       ������������������������       �      �?              @�       ������������������������       ����|���?             &@      S       d                     @�j��e�?u            �f@      T       _                    �?$Q�q�?M            �_@      U       Z                    �?@݈g>h�?.             S@      V       Y                     �?�:�^���?            �F@        W       X                 `��S@�����H�?             2@        ������������������������       �����X�?             @}       ������������������������       �                     &@�       ������������������������       ��>����?             ;@        [       \                    �?��a�n`�?             ?@        ������������������������       �        
             &@        ]       ^                 `f�C@R���Q�?
             4@       ������������������������       ����!pc�?             &@        ������������������������       �                     "@        `       c                    <@p���?             I@        a       b                    7@���N8�?             5@       ������������������������       �        	             0@        ������������������������       �z�G�z�?             @        ������������������������       �                     =@        e       n                    @D7�J��?(            �K@       f       m                 ��Y7@8�A�0��?              F@       g       h                   �"@V������?            �B@        ������������������������       �                      @        i       j                    �?����"�?             =@        ������������������������       �      �?              @        k       l                    .@���N8�?             5@        ������������������������       �      �?              @        ������������������������       �$�q-�?
             *@        ������������������������       �                     @        o       p                    @�C��2(�?             &@        ������������������������       �r�q��?             @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KKqKK��h\�B       0|@     Pp@      n@      O@     �D@      �?      ?@              $@      �?     �h@     �N@      2@       @      @      @      ,@      @     �f@     �J@     `b@      :@     �[@      ,@     �Z@       @      8@      @      @       @      1@      @      @       @      &@      �?     �T@      @     �S@       @      @      �?     �Q@      �?      4@      �?      ,@              @      �?     �I@              @      �?      @      @      B@      (@      &@              9@      (@       @       @      7@      @      .@               @      @      A@      ;@              @      A@      5@      @      @      =@      ,@              @      =@      $@      .@       @      ,@       @      @      @      @       @     `j@     �h@     �e@      K@     �d@      F@     `a@      F@              *@     `a@      ?@      7@      *@       @       @      5@      @      1@      @      (@      @      @              @       @      ]@      2@     @W@      2@      Q@      @     �F@              7@      @      "@       @      ,@      �?      $@              @      �?      9@      .@      @      $@      �?      @      @      @      5@      @      2@      �?       @      �?      $@              @      @      7@              ;@              "@      $@       @      @      @      @      B@      b@       @     �]@      @     @Q@      @     �D@       @      0@       @      @              &@       @      9@      @      <@              &@      @      1@      @       @              "@      �?     �H@      �?      4@              0@      �?      @              =@      <@      ;@      2@      :@      &@      :@               @      &@      2@      @       @      @      0@      @      @      �?      (@      @              $@      �?      @      �?      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��.hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsK}hth)h,K ��h.��R�(KK}��h{�B@         *                 ��%@(����7�?�           @�@      @                           /@�BPԃ�?�             r@       @������������������������       �      �?              @1���                             �?��X)�^�?�            �q@2���                             �?�KM�]�?�            �l@       @                        ���@������?             ;@        ������������������������       �z�G�z�?             $@      @������������������������       ��t����?             1@       @	       
                   �0@�7A��?�             i@      ;@������������������������       �      �?              @      ,@                         ��@<2r�Y�?|             h@       @                          �8@@��8��?!             H@      K@                        ���@���7�?             6@      ?@������������������������       ��C��2(�?             &@      @������������������������       �                     &@      2@������������������������       �                     :@      @                        �1@h�:��T�?[             b@                               ��@���!pc�?             6@                                �=@�8��8��?
             (@      ������������������������       �؇���X�?             @w      ������������������������       �                     @n      ������������������������       �      �?             $@�                                �>@@;�"�?J            �^@                                �4@�g�y��?6            @W@       ������������������������       �r�q��?             2@�      ������������������������       �        *            �R@c                              @3�@r�q��?             >@       ������������������������       ��q�q�?             (@                                �E@�X�<ݺ?             2@      ������������������������       �        
             (@(      ������������������������       �r�q��?             @V              #                   �5@�5��?&             K@       !       "                 ��Y@�C��2(�?             &@       ������������������������       �r�q��?             @A      ������������������������       �                     @�       $       '                  ��@X��ʑ��?            �E@       %       &                  ��@ �o_��?             9@        ������������������������       ����Q��?             @j       ������������������������       �      �?             4@�       (       )                   �>@�<ݚ�?             2@       ������������������������       ��8��8��?	             (@�       ������������������������       �      �?             @�       +       v                    @�-����?           `z@       ,       M                     �?�D&\���?�            �w@        -       0                   �1@�r�K��?c            `d@        .       /                    �?�S����?	             3@        ������������������������       �                      @]       ������������������������       ����!pc�?             &@�       1       B                    �?��E�@�?Z             b@       2       =                 ���S@      �?5            �V@       3       <                    �?p�EG/��?$            �O@       4       ;                   �>@l��
I��?             K@       5       :                   �J@П[;U��?             =@       6       9                 ���=@
;&����?             7@      7       8                   �D@ҳ�wY;�?             1@        ������������������������       �                     @`      ������������������������       ����Q��?             $@:      ������������������������       �                     @;      ������������������������       �r�q��?             @?      ������������������������       �H%u��?             9@I      ������������������������       �                     "@7      >       A                  ޅg@������?             ;@       ?       @                    �?ףp=
�?             4@       ������������������������       �      �?              @!      ������������������������       �                     (@�      ������������������������       �����X�?             @�      C       H                    E@l��
I��?%             K@       D       E                    :@�J�4�?             9@       ������������������������       �և���X�?             @      F       G                    �?�X�<ݺ?             2@       ������������������������       �r�q��?             @,      ������������������������       �                     (@�      I       L                    �?�f7�z�?             =@       J       K                 Ј�U@�q�q�?             2@       ������������������������       �      �?             (@v      ������������������������       �      �?             @�      ������������������������       �                     &@�      N       Y                 `�X.@���=��?�            @k@       O       V                 ��+@���Q��?5            @U@      P       S                    �?������?(            �O@      Q       R                   �3@v�X��?             F@        ������������������������       ����|���?             &@      ������������������������       �"pc�
�?            �@@-      T       U                    :@�}�+r��?             3@       ������������������������       �      �?             @g      ������������������������       �        	             .@�       W       X                    :@��2(&�?             6@        ������������������������       ��z�G��?             $@}       ������������������������       �        	             (@�       Z       u                    @B��仱�?[            �`@       [       \                    !@����1�?W            �_@        ������������������������       �                     .@        ]       r                    �?�f��`��?K            �[@       ^       a                 ��0@������?;            �U@        _       `                 ���/@"pc�
�?	             &@       ������������������������       �؇���X�?             @        ������������������������       �      �?             @        b       g                    �?��=A��?2             S@        c       f                    �?X�<ݚ�?             ;@       d       e                 0��D@և���X�?             5@       ������������������������       ��θ�?             *@        ������������������������       �      �?              @        ������������������������       �                     @        h       o                    �?�J��%�?!            �H@       i       n                    �?�����H�?             ;@       j       m                   �@@@�0�!��?             1@       k       l                    �?���!pc�?
             &@       ������������������������       �����X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     $@        p       q                    �?8�A�0��?             6@       ������������������������       �     ��?             0@        ������������������������       �                     @        s       t                     @      �?             8@        ������������������������       �"pc�
�?             &@        ������������������������       ��	j*D�?             *@        ������������������������       �                     @        w       |                    @������?            �D@       x       {                   �7@��� ��?             ?@       y       z                    �?HP�s��?             9@       ������������������������       �        	             .@        ������������������������       �z�G�z�?             $@        ������������������������       ��q�q�?             @        ������������������������       �                     $@        �t�bh�h)h,K ��h.��R�(KK}KK��h\�B�       �{@      q@     �l@      O@       @      @     @l@      L@     �i@      8@      4@      @       @       @      (@      @      g@      1@      @       @     @f@      .@     �G@      �?      5@      �?      $@      �?      &@              :@             ``@      ,@      0@      @      &@      �?      @      �?      @              @      @     �\@       @     �V@      @      .@      @     �R@              9@      @       @      @      1@      �?      (@              @      �?      6@      @@      �?      $@      �?      @              @      5@      6@      @      2@       @      @      @      .@      ,@      @      &@      �?      @      @     �j@     @j@     �e@     �i@      P@     �X@      @      0@               @      @       @     �N@     �T@     �F@     �F@      C@      9@      C@      0@      0@      *@      &@      (@      &@      @      @              @      @              @      @      �?      6@      @              "@      @      4@       @      2@       @      @              (@      @       @      0@      C@      @      5@      @      @      �?      1@      �?      @              (@      (@      1@      (@      @      "@      @      @      @              &@     �[@     �Z@     �I@      A@      @@      ?@      ?@      *@      @      @      ;@      @      �?      2@      �?      @              .@      3@      @      @      @      (@              N@     @R@     �J@     @R@              .@     �J@      M@     �G@      D@       @      "@      �?      @      �?      @     �F@      ?@      (@      .@      (@      "@      $@      @       @      @              @     �@@      0@      8@      @      ,@      @       @      @      @       @      @      �?      @              $@              "@      *@      "@      @              @      @      2@       @      "@      @      "@      @             �B@      @      ;@      @      7@       @      .@               @       @      @       @      $@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��~hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKkhth)h,K ��h.��R�(KKk��h{�B�         `                 ��gS@l��n�?�           @�@     @       =                    �?�xt��?�           ��@     @                           �?�u�s#�?           {@                                  �;@�1�`jg�?"            �K@        ������������������������       �      �?             ,@      �?                          �=@��P���?            �D@     @                          @@������?             ;@      @������������������������       �@4և���?             ,@      @@	       
                     �?��
ц��?	             *@      6@������������������������       �      �?              @      @������������������������       ����Q��?             @     �i@                          @B@؇���X�?	             ,@      @������������������������       �                      @      0@������������������������       ��q�q�?             @               .                 ��D:@��4k��?�            �w@     @       +                    �?$V�Ap�?�            �q@     @                          �4@(�qEy��?�            Pp@       ������������������������       �                     J@�                                  @�KM�]�?�             j@                                  ?@�U�:��?(            �M@       ������������������������       �                     <@n      ������������������������       ��חF�P�?             ?@�                                �;@��cˣ��?b            �b@                                 �7@d}h���?             E@       ������������������������       ��C��2(�?             6@�                              ��L@��Q��?             4@       ������������������������       ��q�q�?             "@      ������������������������       ��C��2(�?             &@                               s�@�>����?F             [@       ������������������������       �                     7@(             "                 �Y5@��O���?8            @U@               !                 ��@      �?             0@      ������������������������       ����!pc�?             &@3      ������������������������       �z�G�z�?             @A      #       $                   �<@p��%���?-            @Q@        ������������������������       �                     B@�       %       &                 @3�@<���D�?            �@@        ������������������������       ��<ݚ�?             "@j       '       *                 ���"@�8��8��?             8@       (       )                   �@@�}�+r��?             3@        ������������������������       �؇���X�?             @�       ������������������������       �                     (@�       ������������������������       �z�G�z�?             @$       ,       -                    )@���Q��?             9@        ������������������������       ��C��2(�?             &@       ������������������������       �                     ,@-       /       8                     �?���j��?9             W@       0       5                   �>@Fx$(�?              I@       1       4                   �J@X�<ݚ�?             ;@       2       3                 `f�;@�d�����?             3@       ������������������������       �ףp=
�?             $@�       ������������������������       �X�<ݚ�?             "@�       ������������������������       �      �?              @�       6       7                    �?�㙢�c�?             7@       ������������������������       �                     (@�       ������������������������       ����|���?             &@`      9       <                   �C@r�q��?             E@       :       ;                    +@�E��ӭ�?             2@      ������������������������       ��eP*L��?             &@?      ������������������������       �                     @I      ������������������������       ��8��8��?             8@7      >       G                     @ �
��?~            �i@        ?       B                     �?�zvܰ?9             V@       @       A                  �>I@@4և���?             <@       ������������������������       ��q�q�?             @�      ������������������������       �                     6@�      C       F                   �;@ �.�?Ƞ?(             N@        D       E                    �?���7�?             6@       ������������������������       �      �?              @      ������������������������       �        	             ,@-      ������������������������       �                     C@,      H       [                    �?z4��f��?E            @]@      I       X                   �<@�q�Q�?7             X@       J       W                 �16@|�U&k�?,            �R@       K       P                   �8@���!pc�?(            �P@       L       O                   �4@�J�4�?             9@      M       N                    �?�	j*D�?
             *@       ������������������������       ����Q��?             @�      ������������������������       �      �?              @�      ������������������������       �                     (@�      Q       V                    �?#z�i��?            �D@       R       U                    �?�t����?             A@      S       T                    �?��<b���?             7@      ������������������������       �������?	             1@%      ������������������������       �r�q��?             @g      ������������������������       ��eP*L��?             &@�       ������������������������       �և���X�?             @y       ������������������������       �      �?              @}       Y       Z                    @"pc�
�?             6@       ������������������������       �����X�?             ,@        ������������������������       �                      @        \       _                    7@؇���X�?             5@       ]       ^                 `f�=@�C��2(�?	             &@       ������������������������       �                     @        ������������������������       �z�G�z�?             @        ������������������������       �z�G�z�?             $@        a       f                    �?�MI8d�?-            �R@        b       e                    �?D�n�3�?             3@       c       d                 �U�X@X�Cc�?	             ,@        ������������������������       �      �?             @        ������������������������       �      �?              @        ������������������������       ����Q��?             @        g       h                  "�b@ �Jj�G�?             �K@       ������������������������       �                    �C@        i       j                 `D�g@      �?
             0@        ������������������������       �r�q��?             @        ������������������������       �                     $@        �t�bh�h)h,K ��h.��R�(KKkKK��h\�B�       {@     pq@     Pz@      k@     pv@     �R@     �C@      0@      @      @      @@      "@      4@      @      *@      �?      @      @      @      @      @       @      (@       @       @              @       @      t@      M@     �o@      @@     �m@      6@      J@             `g@      6@      K@      @      <@              :@      @     �`@      1@     �@@      "@      4@       @      *@      @      @      @      $@      �?      Y@       @      7@             @S@       @      (@      @       @      @      @      �?     @P@      @      B@              =@      @      @       @      6@       @      2@      �?      @      �?      (@              @      �?      .@      $@      �?      $@      ,@             �P@      :@      ?@      3@      (@      .@      @      ,@      �?      "@      @      @      @      �?      3@      @      (@              @      @     �A@      @      *@      @      @      @      @              6@       @      O@     �a@      @     @U@       @      :@       @      @              6@      �?     �M@      �?      5@      �?      @              ,@              C@     �M@      M@     �D@     �K@      7@     �I@      2@      H@      @      5@      @      "@      @       @      �?      @              (@      ,@      ;@      $@      8@      @      2@      @      *@      �?      @      @      @      @      @      @      @      2@      @      $@      @       @              2@      @      $@      �?      @              @      �?       @       @      (@      O@      &@       @      "@      @      @      @      @       @       @      @      �?      K@             �C@      �?      .@      �?      @              $@�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��.hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKwhth)h,K ��h.��R�(KKw��h{�B�         *                     @<��z��?�           @�@                                   �?
;&����?�             t@DԤ�                             $@�-���?             i@        ������������������������       �                     (@      �?                            �?��[�p�?y            �g@      @                          �K@��|�	��?<            �V@     "@                           �?�4F����?5            �T@      �?                           �?|��?���?             ;@     @	       
                 `f�C@և���X�?             5@        ������������������������       ����!pc�?             &@      �?                          �?@���Q��?             $@      $@������������������������       ����Q��?             @      3@������������������������       ����Q��?             @      @������������������������       ��q�q�?             @      @                           >@�rF���?#            �K@        ������������������������       ������?             5@      :@                           �?�t����?             A@      ������������������������       �z�G�z�?             4@�      ������������������������       �և���X�?	             ,@�      ������������������������       �X�<ݚ�?             "@w                                 �?�$��y��?=            @X@                                �I@      �?,             R@                                @A@\#r��?'            �N@                                �;@��E�B��?            �G@      ������������������������       �`Jj��?             ?@�                                 @      �?             0@       ������������������������       �                     @      ������������������������       ����|���?             &@      ������������������������       �        
             ,@�      ������������������������       ����!pc�?             &@(      ������������������������       �                     9@V              %                     �?�.ߴ#�?S            �^@      !       "                    �?$�q-�?*            @P@      ������������������������       �        !             I@A      #       $                   �7@�q�q�?	             .@        ������������������������       �      �?             @�       ������������������������       ��<ݚ�?             "@v       &       )                   �*@0�)AU��?)            �L@        '       (                   �;@@4և���?             ,@        ������������������������       �      �?             @�       ������������������������       �        	             $@�       ������������������������       �                    �E@�       +       v                   �C@r9��X��?�            `x@       ,       _                    �?b��A���?�            �v@       -       N                   �;@L�{[��?�            �n@       .       M                    �?��n��?T            @_@       /       L                    �?�ψX�F�?N            @\@       0       G                 ��i%@~	~���?G            �X@       1       F                 ��Y @�?a/��?;            �T@       2       A                   �8@��R[s�?1            �Q@       3       4                    �?�rF���?%            �K@        ������������������������       ����Q��?             @�       5       >                   �5@j�q����?!             I@       6       ;                   �3@�<ݚ�?             B@      7       8                   �1@R���Q�?             4@        ������������������������       ��<ݚ�?             "@`      9       :                   �@�C��2(�?
             &@      ������������������������       �                     @;      ������������������������       �      �?             @?      <       =                   �4@     ��?
             0@       ������������������������       �և���X�?             @7      ������������������������       ��<ݚ�?             "@G       ?       @                 p�@@4և���?	             ,@       ������������������������       �؇���X�?             @!      ������������������������       �                     @�      B       E                 ��L@���Q��?             .@      C       D                 ���@�eP*L��?             &@        ������������������������       �      �?             @8      ������������������������       ����Q��?             @      ������������������������       �                     @-      ������������������������       �        
             *@,      H       I                    ,@���Q��?             .@       ������������������������       �                     @�       J       K                 03�0@�q�q�?             "@        ������������������������       �z�G�z�?             @v      ������������������������       �      �?             @�      ������������������������       �                     .@�      ������������������������       �                     (@�      O       \                   �>@Xny��?R            �^@      P       [                 03�6@���1j	�?9            �U@      Q       T                    �?P���Q�?4             T@        R       S                   @@�����H�?             2@      ������������������������       ��8��8��?	             (@-      ������������������������       �r�q��?             @%      U       V                  sW@�g�y��?'             O@       ������������������������       ��C��2(�?             &@�       W       X                 ��) @���J��?            �I@       ������������������������       �                    �@@}       Y       Z                    �?�X�<ݺ?             2@       ������������������������       �$�q-�?             *@        ������������������������       �                     @        ������������������������       �r�q��?             @        ]       ^                   @@@      �?             B@        ������������������������       ��q�q�?
             (@        ������������������������       ��8��8��?             8@        `       e                 �̌@~}e}b �?D            �\@        a       b                   �5@R�}e�.�?             :@        ������������������������       �X�<ݚ�?             "@        c       d                 ���@@�0�!��?             1@        ������������������������       �                     @        ������������������������       ��z�G��?             $@        f       s                 ��Y7@�VM�?3            @V@       g       n                 ��.@4�.�A�?&            �O@       h       i                    3@�θ�?            �C@        ������������������������       ��eP*L��?             &@        j       m                 P��%@ �Cc}�?             <@       k       l                 @3�@P���Q�?
             4@        ������������������������       �r�q��?             @        ������������������������       �                     ,@        ������������������������       �      �?              @        o       r                    �?�q�q�?             8@       p       q                    �?      �?
             0@        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �      �?              @        t       u                 ��T?@ȵHPS!�?             :@       ������������������������       �                     1@        ������������������������       ��q�q�?             "@        ������������������������       �                     <@        �t�bh�h)��     h,K ��h.��R�(KKwKK��h\�Bp       p|@     p@     @c@      e@     �b@      J@              (@     �b@      D@      N@      ?@      L@      :@      *@      ,@      "@      (@      @       @      @      @      @       @      @       @      @       @     �E@      (@      3@       @      8@      $@      0@      @       @      @      @      @      V@      "@     �O@      "@     �K@      @     �D@      @      =@       @      (@      @      @              @      @      ,@               @      @      9@              @      ]@      @      N@              I@      @      $@      @      @       @      @      �?      L@      �?      *@      �?      @              $@             �E@     �r@     @V@     q@     @V@     �i@     �D@     �X@      ;@     �U@      ;@     �Q@      ;@     @P@      2@      J@      2@     �E@      (@       @      @     �D@      "@      <@       @      1@      @      @       @      $@      �?      @              @      �?      &@      @      @      @      @       @      *@      �?      @      �?      @              "@      @      @      @      @      @       @      @      @              *@              @      "@              @      @      @      @      �?       @       @      .@              (@              [@      ,@     @T@      @      S@      @      0@       @      &@      �?      @      �?      N@       @      $@      �?      I@      �?     �@@              1@      �?      (@      �?      @              @      �?      ;@      "@      @      @      6@       @     �P@      H@      @      3@      @      @      @      ,@              @      @      @      N@      =@     �B@      :@      >@      "@      @      @      9@      @      3@      �?      @      �?      ,@              @       @      @      1@      @      (@               @      @      @      @      @      7@      @      1@              @      @      <@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�DhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKmhth)h,K ��h.��R�(KKm��h{�B@         `                 �U�R@��6���?�           @�@              #                     @8kT���?�           ��@      @                           �?(ǯt��?�            �k@      @                           1@��Hg���?Z            �`@      @������������������������       �      �?              @      @                           �?@w��_m�?V            �_@     @                          �:@      �?N             [@      @������������������������       �      �?             8@      ]@	                            �?����X�?=             U@     @
                           �?�n_Y�K�?%             J@      @������������������������       ��z�G��?             $@     @V@                           �?�D����?             E@     ;@                          �J@�Gi����?            �B@     @                          �>@     ��?             @@      @                          �9@      �?             8@      @������������������������       �                     @      �?                          �E@r�q��?
             2@       ������������������������       �                     $@�      ������������������������       �      �?              @�      ������������������������       �                      @w      ������������������������       �                     @n      ������������������������       ����Q��?             @�                                �<@      �?             @@       ������������������������       �      �?             (@�                                �@@P���Q�?             4@       ������������������������       �                     "@c                                �B@�C��2(�?
             &@       ������������������������       �      �?             @      ������������������������       �                     @�      ������������������������       �                     3@(             "                   �;@XB���?9            �U@               !                    6@�#-���?            �A@       ������������������������       ��q�q�?             "@3      ������������������������       �                     :@A      ������������������������       �        "             J@�       $       )                    @S�o��?�            py@        %       (                 @3�4@��X��?             <@       &       '                    �?ףp=
�?
             4@        ������������������������       �                     "@�       ������������������������       �"pc�
�?             &@�       ������������������������       �      �?              @�       *       K                    �?��}�v��?�            �w@       +       H                 �T�I@�θV�?�            @q@       ,       G                   @@@8�B�n�?�            pp@       -       F                   �?@$�q-�?~             j@       .       ;                   �;@�����?x            �h@       /       :                   �9@L紂P�?>            �Y@       0       5                 ��@�q��/��?7             W@        1       2                   �5@Pa�	�?            �@@        ������������������������       �                     *@�       3       4                 �Y�@P���Q�?
             4@        ������������������������       �r�q��?             @�       ������������������������       �                     ,@�       6       9                    0@@�r-��?&            �M@      7       8                   �5@d}h���?             E@       ������������������������       �r֛w���?             ?@`      ������������������������       ��C��2(�?             &@:      ������������������������       �        	             1@;      ������������������������       ����Q��?             $@?      <       =                    �?h�a��?:            @X@       ������������������������       �                    �A@7      >       E                    �?6uH���?!             O@       ?       D                   @<@�C��2(�?            �K@      @       C                 pf� @�����?             E@      A       B                 �?�@�r����?             >@      ������������������������       �      �?	             0@�      ������������������������       �؇���X�?             ,@8       ������������������������       �                     (@8      ������������������������       �$�q-�?             *@      ������������������������       �                     @-      ������������������������       �X�<ݚ�?             "@,      ������������������������       �        $            �K@�      I       J                    �?�n_Y�K�?	             *@       ������������������������       �r�q��?             @�       ������������������������       �                     @v      L       M                   �-@D;����?C            �Y@       ������������������������       ������H�?             "@�      N       [                    �?��V�I��?=            �W@      O       P                    �?p�EG/��?)            �O@       ������������������������       �X�<ݚ�?             "@�      Q       Z                    �?��}*_��?"             K@       R       S                   �4@r�qG�?             H@       ������������������������       ��eP*L��?             &@-      T       U                    �?V������?            �B@       ������������������������       �     ��?             0@g      V       W                   �@�ՙ/�?             5@        ������������������������       �                     $@y       X       Y                   �;@���!pc�?             &@        ������������������������       �z�G�z�?             @�       ������������������������       ��q�q�?             @        ������������������������       �      �?             @        \       ]                    �?`՟�G��?             ?@        ������������������������       ��q�q�?             (@        ^       _                  ��8@p�ݯ��?             3@        ������������������������       ��<ݚ�?             "@        ������������������������       �                     $@        a       f                    �?��Lɿ��?1            �T@       b       e                 0w�a@���N8�?             E@       c       d                    �?ףp=
�?             4@        ������������������������       �      �?              @        ������������������������       �        	             (@        ������������������������       �                     6@        g       l                   �H@��r._�?            �D@       h       k                    �?      �?             @@        i       j                 pޅV@X�<ݚ�?             "@        ������������������������       ����Q��?             @        ������������������������       �      �?             @        ������������������������       �                     7@        ������������������������       ��q�q�?             "@        �t�bh�h)h,K ��h.��R�(KKmKK��h\�B�       Pz@     0r@     �y@      k@     @Z@     @]@     �Y@     �@@       @      @      Y@      ;@     @T@      ;@      5@      @      N@      8@      @@      4@      @      @      9@      1@      6@      .@      1@      .@      "@      .@      @              @      .@              $@      @      @       @              @              @       @      <@      @      "@      @      3@      �?      "@              $@      �?      @      �?      @              3@              @      U@      @      @@      @      @              :@              J@     0s@      Y@      "@      3@       @      2@              "@       @      "@      @      �?     �r@     @T@      o@      <@      n@      7@      g@      7@     �f@      3@      V@      ,@     �T@      $@      @@      �?      *@              3@      �?      @      �?      ,@              I@      "@     �@@      "@      7@       @      $@      �?      1@              @      @      W@      @     �A@             �L@      @      I@      @      C@      @      :@      @      ,@       @      (@       @      (@              (@      �?      @              @      @     �K@               @      @      �?      @      @              I@     �J@       @      �?      E@      J@      9@      C@      @      @      4@      A@      1@      ?@      @      @      &@      :@      @      *@       @      *@              $@       @      @      @      �?      @       @      @      @      1@      ,@      @      @      (@      @       @      @      $@              "@     �R@       @      D@       @      2@       @      @              (@              6@      @      A@      @      <@      @      @       @      @       @       @              7@      @      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ���MhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKshth)h,K ��h.��R�(KKs��h{�B�         2                     @�U��h��?�           @�@                                  �1@�n�q�Z�?�            `s@                                   �?��a�n`�?             ?@     �U@������������������������       ��q�q�?             @      6@                            �?`2U0*��?             9@        ������������������������       �؇���X�?             @      @������������������������       �                     2@      �?       %                    �?����?�            pq@     @@	                           �?z�G�z�?k             d@     Y@
                           �?��j���?O            �[@     "@                        ���<@r�q��?H            �Y@     7@                          �@@�S(��d�?4            @S@     $@                            �?��Y��]�?            �D@      �?������������������������       �                     $@       @                           5@�g�y��?             ?@      @������������������������       �      �?              @      @������������������������       �                     7@Z                                �E@4?,R��?             B@                                 �B@�q�q�?
             .@       ������������������������       �      �?              @w      ������������������������       �����X�?             @n      ������������������������       �                     5@�                                 @@� �	��?             9@                                 @>@�q�q�?	             (@       ������������������������       �      �?             @�      ������������������������       �r�q��?             @c                                �@@�θ�?             *@      ������������������������       �؇���X�?             @      ������������������������       ��q�q�?             @�      ������������������������       �                     "@(             $                     �?~���L0�?            �H@              #                   �G@l��[B��?             =@      !       "                   �;@�ՙ/�?             5@       ������������������������       �؇���X�?             @A      ������������������������       �؇���X�?             ,@�       ������������������������       �      �?              @�       ������������������������       �                     4@v       &       /                   �H@ ����?N            �]@       '       (                    �?@��!�Q�?B            @Z@       ������������������������       �        #             L@�       )       .                    �?@�E�x�?            �H@       *       +                     �?h�����?             <@       ������������������������       �                     1@$       ,       -                   �;@�C��2(�?             &@        ������������������������       �r�q��?             @       ������������������������       �                     @-       ������������������������       �                     5@]       0       1                   @I@@4և���?             ,@        ������������������������       �      �?             @A       ������������������������       �                     $@�       3       j                    �?!��)��?�             y@       4       ;                   �0@h���e0�?�             v@        5       8                    �?8^s]e�?             =@        6       7                 `f�@�r����?	             .@       ������������������������       �r�q��?             @�       ������������������������       ������H�?             "@`      9       :                    �?      �?
             ,@       ������������������������       �z�G�z�?             @;      ������������������������       ��q�q�?             "@?      <       ]                 `�X.@$�	W��?�            0t@      =       V                    �?RB)��.�?�             p@      >       S                   @@@hD=�$��?�            �i@       ?       R                 pF�'@��r._�?g            �d@      @       O                   �<@��ۭ���?b            �c@      A       F                 �Y�@�Ra����?S            �`@       B       C                    7@      �?             4@       ������������������������       �؇���X�?             @8       D       E                 ���@�	j*D�?
             *@       ������������������������       ��q�q�?             @      ������������������������       �����X�?             @-      G       N                    �?4և����?E             \@      H       I                   �:@�NW���?A            �Z@      ������������������������       � =[y��?%             Q@�       J       K                    �?�?�'�@�?             C@        ������������������������       �                     "@v      L       M                 ��) @д>��C�?             =@      ������������������������       �                     6@�      ������������������������       �����X�?             @�      ������������������������       ��q�q�?             @�      P       Q                   �?@�q�����?             9@      ������������������������       ���.k���?	             1@�       ������������������������       �      �?              @      ������������������������       �                     @-      T       U                 �?�@�Ń��̧?             E@      ������������������������       �                     :@g      ������������������������       �      �?             0@�       W       \                 �̌@��B����?"             J@        X       Y                 ���@ �o_��?             9@        ������������������������       �                      @�       Z       [                    �?j���� �?
             1@        ������������������������       �؇���X�?             @        ������������������������       ����Q��?             $@        ������������������������       �������?             ;@        ^       e                    �?�G\�c�?&            @P@       _       d                    �?�<ݚ�?             B@       `       c                    �?R�}e�.�?             :@       a       b                 �T)D@��
ц��?             *@        ������������������������       �z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     *@        ������������������������       �ףp=
�?             $@        f       g                    �?J�8���?             =@        ������������������������       �     ��?	             0@        h       i                    �?��
ц��?	             *@       ������������������������       �؇���X�?             @        ������������������������       �                     @        k       n                 03�7@ "��u�?             I@        l       m                    7@"pc�
�?             &@        ������������������������       �      �?             @        ������������������������       �؇���X�?             @        o       r                 ��p@@ ���J��?            �C@        p       q                    @�}�+r��?             3@        ������������������������       �      �?              @        ������������������������       �                     &@        ������������������������       �                     4@        �t�bh�h)h,K ��h.��R�(KKsKK��h\�B0       �z@     �q@     �`@      f@      @      <@       @      @      �?      8@      �?      @              2@     @`@     �b@      `@      @@     �W@      1@     @U@      1@     �Q@      @      D@      �?      $@              >@      �?      @      �?      7@              ?@      @      $@      @      @      @      @       @      5@              ,@      &@      @       @      @      @      �?      @      $@      @      @      �?      @       @      "@              A@      .@      ,@      .@      *@       @      �?      @      (@       @      �?      @      4@               @     @]@      �?      Z@              L@      �?      H@      �?      ;@              1@      �?      $@      �?      @              @              5@      �?      *@      �?      @              $@     �r@      Z@     `o@     @Y@      "@      4@       @      *@      �?      @      �?       @      @      @      @      �?      @      @     @n@     @T@     �i@      K@      f@      =@      a@      <@      `@      <@     @]@      .@      .@      @      @      �?      "@      @      @       @      @       @     �Y@      $@     �X@       @     @P@      @     �@@      @      "@              8@      @      6@               @      @      @       @      (@      *@      "@       @      @      @      @             �D@      �?      :@              .@      �?      ;@      9@      @      2@               @      @      $@      �?      @      @      @      4@      @      C@      ;@      <@       @      3@      @      @      @      @      �?       @      @      *@              "@      �?      $@      3@      @      *@      @      @      �?      @      @             �G@      @      "@       @      @      �?      @      �?      C@      �?      2@      �?      @      �?      &@              4@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ9M�hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKmhth)h,K ��h.��R�(KKm��h{�B@         B                    �?���y�?�           @�@              +                 ��$:@�r�5S��?*            }@    �b@                           $@PU�k ��?�            0t@     �@@������������������������       �                     &@      9@       *                    �?��-�=��?�            �s@     @       	                    �?Y��!�?�             r@       @                           ;@z�G�z�?            �A@      �?������������������������       ����Q��?             $@      .@������������������������       �H%u��?             9@      @
                            �?`�H�/��?�            �o@      L@������������������������       �                     @      $@       '                   �*@��I�?�             o@     *@                        �?�@\�����?�            @j@     @Y@                          @@@�c:��?@             W@      @                            @h��@D��?1            �Q@     @T@������������������������       �                     @      <@                           �?     ��?-             P@       ������������������������       �      �?
             0@�                              �{@      �?#             H@                                �8@     ��?             @@                              �?$@���N8�?             5@      ������������������������       �        	             *@�      ������������������������       �      �?              @�      ������������������������       ��eP*L��?             &@�      ������������������������       �                     0@�      ������������������������       �                     5@c                                �1@(2��R�?K            �]@       ������������������������       ����Q��?             @                               @3�@4��Q���?G            @\@                                 @A@�q�q�?	             (@      ������������������������       �����X�?             @V      ������������������������       ����Q��?             @J      !       "                     @��T�u��?>            @Y@       ������������������������       �*
;&���?             G@A      #       $                 @Q!@h㱪��?#            �K@       ������������������������       �                     @@�       %       &                 ���!@���}<S�?             7@        ������������������������       �"pc�
�?             &@j       ������������������������       �                     (@�       (       )                 03�6@�7��?            �C@       ������������������������       �                     ;@�       ������������������������       �r�q��?             (@�       ������������������������       �                     6@$       ,       ;                    �?$�}�$>�?W            �a@       -       :                     @k�q��?6            @U@       .       3                   �>@�;u�,a�?1            �S@        /       2                  I>@��Zy�?            �C@       0       1                 `f�:@     ��?             @@        ������������������������       �ҳ�wY;�?	             1@A       ������������������������       �������?
             .@�       ������������������������       �                     @�       4       7                    �?�z�G��?             D@       5       6                 `fS@�8��8��?             8@       ������������������������       �                     .@      ������������������������       ��<ݚ�?             "@�       8       9                    �?      �?             0@       ������������������������       �      �?              @:      ������������������������       �      �?              @;      ������������������������       �r�q��?             @?      <       A                     @\-��p�?!             M@       =       >                    �?�	j*D�?             :@       ������������������������       �և���X�?             @G       ?       @                     �?���y4F�?             3@      ������������������������       �"pc�
�?             &@!      ������������������������       �      �?              @�      ������������������������       �                     @@�      C       d                    �? ͵H��?�            �n@       D       _                 ��	6@�L���?v             h@      E       J                     @b�2�tk�?G            �_@       F       I                   �*@��a�n`�?             ?@      G       H                 `f�)@���7�?             6@       ������������������������       �                     (@�      ������������������������       �ףp=
�?             $@�       ������������������������       ��<ݚ�?             "@�       K       \                    �?��C����?7            �W@      L       Y                    .@bf@����?,            �S@      M       X                    �?�\����?$            �P@      N       Q                  s�@l`N���?            �J@       O       P                 03s@؇���X�?	             ,@       ������������������������       �z�G�z�?             @�      ������������������������       ������H�?             "@�       R       S                    �?Hث3���?            �C@       ������������������������       �      �?             ,@-      T       W                   �;@�q�����?             9@      U       V                 pf� @      �?	             0@      ������������������������       ��z�G��?             $@�       ������������������������       �      �?             @y       ������������������������       ��<ݚ�?             "@}       ������������������������       �                     *@�       Z       [                 @3�/@$�q-�?             *@        ������������������������       �                     @        ������������������������       �؇���X�?             @        ]       ^                 @�+@      �?             0@       ������������������������       ��q�q�?             "@        ������������������������       �                     @        `       c                 ��A@0�,���?/            �P@        a       b                    �?      �?             0@       ������������������������       �z�G�z�?             $@        ������������������������       �                     @        ������������������������       �        "            �I@        e       f                    �?��k��?!            �J@        ������������������������       �                     @        g       h                 03�;@�q�q��?             H@        ������������������������       ��8��8��?             (@        i       j                    )@�<ݚ�?             B@        ������������������������       �      �?             0@        k       l                 ���Q@��Q��?             4@       ������������������������       �$�q-�?             *@        ������������������������       �؇���X�?             @        �t�bh�h)h,K ��h.��R�(KKmKK��h\�B�       �|@      p@     �w@     �V@     �q@     �E@              &@     �q@      @@      p@      @@      <@      @      @      @      6@      @     �l@      9@      @              l@      9@     `g@      7@     @U@      @      P@      @      @             �L@      @      .@      �?      E@      @      :@      @      4@      �?      *@              @      �?      @      @      0@              5@             �Y@      0@      @       @     �X@      ,@      @      @      @       @       @      @      W@      "@     �C@      @     �J@       @      @@              5@       @      "@       @      (@             �B@       @      ;@              $@       @      6@              X@     �G@      G@     �C@     �F@      A@      1@      6@      1@      .@      @      &@      &@      @              @      <@      (@      6@       @      .@              @       @      @      $@       @      @      @      @      �?      @      I@       @      2@       @      @      @      .@      @      "@       @      @       @      @@              T@     �d@     �I@     �a@     �H@     @S@      @      <@      �?      5@              (@      �?      "@       @      @      G@     �H@      B@     �E@     �A@      ?@      6@      ?@       @      (@      �?      @      �?       @      4@      3@      @      @      *@      (@      @      $@      @      @      @      @      @       @      *@              �?      (@              @      �?      @      $@      @      @      @      @               @     @P@       @      ,@       @       @              @             �I@      =@      8@              @      =@      3@      �?      &@      <@       @      .@      �?      *@      @      (@      �?      �?      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJpVhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKqhth)h,K ��h.��R�(KKq��h{�B@         N                    �?T�����?�           @�@                                  !@���B�?,           p~@     �S@                           �?r٣����?            �@@        ������������������������       ��q�q�?             "@                                   �?�8��8��?             8@     @������������������������       �        
             3@      @������������������������       ����Q��?             @       @       9                 ��D:@8R����?           `|@     @	       ,                 �&@@Iu]���?�            �u@       
                            �?`7nev^�?�            @p@       @������������������������       �                     $@     �G@                          �0@��f�R@�?�            @o@      .@������������������������       ��z�G��?             $@      (@                           �?2Tv���?�             n@      $@                        ���@��<b���?             7@       @������������������������       �����X�?             @       @������������������������       �     ��?	             0@Z                               ��@��a�n`�?�             k@                                  �?`�q�0ܴ?            �G@       ������������������������       �                     @w                                �;@������?            �D@                                  7@�����?             5@      ������������������������       �                     0@�      ������������������������       ����Q��?             @�      ������������������������       �                     4@�             +                    �?<���i�?f            @e@                                 �<@�Uk���?a            �d@                                @@�q-�?:             Z@                                  �?�S����?             3@      ������������������������       ��C��2(�?             &@(      ������������������������       �      �?              @V      ������������������������       �Pq�����?-            @U@J      !       "                    �?��.��?'            �N@       ������������������������       �؇���X�?             @A      #       &                   @@@r�q��?"             K@        $       %                 @3�@��Q��?             4@        ������������������������       �      �?              @v       ������������������������       �r�q��?             (@j       '       *                   �J@�IєX�?             A@       (       )                   @C@XB���?             =@       ������������������������       �        	             .@�       ������������������������       �@4և���?             ,@�       ������������������������       �z�G�z�?             @$       ������������������������       ����Q��?             @       -       2                   �?@ p�/��?>            @V@       .       /                  �v6@@3����?%             K@       ������������������������       �                     E@]       0       1                  ��8@�8��8��?	             (@       ������������������������       �      �?              @A       ������������������������       �                     @�       3       6                   �*@�#-���?            �A@        4       5                   �F@r�q��?	             (@       ������������������������       ����Q��?             @�       ������������������������       �                     @      7       8                 03�9@�nkK�?             7@       ������������������������       �                     0@`      ������������������������       �؇���X�?             @:      :       =                    :@n�����?>            @Z@       ;       <                    �?�r����?
             .@       ������������������������       �����X�?             @I      ������������������������       �                      @7      >       E                    @@���Q��?4            �V@        ?       @                    �?��Zy�?            �C@       ������������������������       �                     @!      A       D                     �?     ��?             @@      B       C                   �>@      �?	             4@       ������������������������       �ףp=
�?             $@8       ������������������������       ����Q��?             $@8      ������������������������       ��q�q�?             (@      F       M                    �?t�F�}�?             �I@      G       J                   �G@V������?            �B@       H       I                  I=@ףp=
�?
             4@       ������������������������       �      �?              @�       ������������������������       �                     (@�       K       L                    K@��.k���?             1@      ������������������������       ����!pc�?             &@�      ������������������������       �r�q��?             @�      ������������������������       �d}h���?             ,@�      O       j                   �=@������?�             l@      P       [                     @nM`����?\            @a@       Q       T                    6@ܷ��?��?'             M@        R       S                 `f�)@      �?             0@       ������������������������       �                     @-      ������������������������       ����Q��?             $@%      U       V                    �?���N8�?             E@       ������������������������       �        
             2@�       W       X                    �?�8��8��?             8@        ������������������������       �                     @}       Y       Z                 ���`@�����H�?             2@       ������������������������       �        
             ,@        ������������������������       �      �?             @        \       _                  ��@     ��?5             T@        ]       ^                    4@��<b���?             7@        ������������������������       �      �?              @        ������������������������       ���S�ۿ?
             .@        `       a                    @��U/��?'            �L@        ������������������������       ��<ݚ�?             "@        b       e                   �:@�q�q�?             H@       c       d                    �?$�q-�?             :@        ������������������������       ��<ݚ�?             "@        ������������������������       �                     1@        f       g                    �?���|���?             6@        ������������������������       ����Q��?             $@        h       i                     @�q�q�?	             (@       ������������������������       ��q�q�?             @        ������������������������       �                     @        k       n                   @C@ܷ��?��?4            �U@        l       m                 `ff.@`Ql�R�?            �G@        ������������������������       ������H�?             "@        ������������������������       �                     C@        o       p                     @z�G�z�?             D@       ������������������������       �                     ?@        ������������������������       ������H�?             "@        �t�bh�h)h,K ��h.��R�(KKqKK��h\�B       0|@     Pp@     px@      X@       @      9@      @      @       @      6@              3@       @      @     �w@     �Q@     �s@     �@@     �l@      =@      $@             �k@      =@      @      @     �j@      :@      2@      @      @       @      *@      @     �h@      5@     �F@       @      @             �C@       @      3@       @      0@              @       @      4@             �b@      3@     �b@      1@     @X@      @      0@      @      $@      �?      @       @     @T@      @     �I@      $@      @      �?     �F@      "@      *@      @      @      @      $@       @      @@       @      <@      �?      .@              *@      �?      @      �?      @       @     @U@      @     �J@      �?      E@              &@      �?      @      �?      @              @@      @      $@       @      @       @      @              6@      �?      0@              @      �?     �P@      C@      *@       @      @       @       @              K@      B@      1@      6@      @              $@      6@      @      .@      �?      "@      @      @      @      @     �B@      ,@      :@      &@      2@       @      @       @      (@               @      "@      @       @      @      �?      &@      @      N@     �d@     �I@     �U@      @      J@      @      (@              @      @      @       @      D@              2@       @      6@              @       @      0@              ,@       @       @     �F@     �A@      @      2@      @      @      �?      ,@      D@      1@       @      @      C@      $@      8@       @      @       @      1@              ,@       @      @      @       @      @       @      @      @              "@     �S@      �?      G@      �?       @              C@       @      @@              ?@       @      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKchth)h,K ��h.��R�(KKc��h{�B�         $                  �#@T�����?�           @�@                                   �?X�.;v��?�            �q@      @                          �=@.}Z*�?/            �Q@�y��                             1@�p����?)            �N@ #y��  ������������������������       ��<ݚ�?             "@                                   �?�n_Y�K�?$             J@      @                          �7@�r����?             >@      @������������������������       �      �?             @      @	       
                    �?ȵHPS!�?             :@      @������������������������       �ףp=
�?	             $@      �?������������������������       �      �?             0@       @������������������������       ����!pc�?             6@      �?������������������������       �                     $@       @                           �?�8a$M��?�            �j@                                 �8@l�oA�?r            �f@       @                        ��Y @����˵�?#            �M@                               @3�@�˹�m��?             C@                                �4@h�����?             <@       ������������������������       �        	             *@�                               s@��S�ۿ?
             .@       ������������������������       �                     @n      ������������������������       �      �?              @�      ������������������������       �z�G�z�?             $@�      ������������������������       �                     5@�                                �;@f>�cQ�?O            �^@                               ��]@�ՙ/�?             5@       ������������������������       �      �?             (@      ������������������������       ��<ݚ�?             "@                                  @ܴD��?A            @Y@       ������������������������       �                     &@(      ������������������������       ������H�?:            �V@V              #                   �"@:ɨ��?            �@@      !       "                   �;@�û��|�?             7@      ������������������������       �      �?	             0@A      ������������������������       �؇���X�?             @�       ������������������������       �ףp=
�?             $@�       %       L                     @x>ԛ/��?	           �z@       &       /                   �,@r�q��?�             r@        '       ,                    �?�q�q�?#             N@       (       )                    &@؇���X�?             E@        ������������������������       ��q�q�?             "@�       *       +                    =@�C��2(�?            �@@        ������������������������       �d}h���?	             ,@$       ������������������������       �        	             3@       -       .                    :@�<ݚ�?             2@        ������������������������       �      �?              @-       ������������������������       �                     $@]       0       G                    �?��#Zv�?�            �l@       1       2                   �3@���W9�?S            ``@        ������������������������       �z�G�z�?             $@�       3       F                  D�_@*AA,�P�?N            @^@       4       C                 Ј�U@�/e�U��?I            �[@       5       >                     �?���|�?A            @X@       6       =                    �?@i��M��?+            @P@      7       8                    @@Z�K�D��?             �G@       ������������������������       �� �	��?             9@`      9       <                 �UP@��2(&�?             6@      :       ;                 ���D@$�q-�?             *@       ������������������������       �r�q��?             @?      ������������������������       �                     @I      ������������������������       ��<ݚ�?             "@7      ������������������������       ��<ݚ�?             2@G       ?       B                    @@      �?             @@       @       A                    �?      �?             0@      ������������������������       ��<ݚ�?             "@�      ������������������������       �����X�?             @�      ������������������������       �                     0@8       D       E                   �B@����X�?             ,@       ������������������������       �z�G�z�?             $@      ������������������������       �      �?             @-      ������������������������       �                     $@,      H       I                    �?�a�O�?9            @X@      ������������������������       �        0            @T@�       J       K                   �W@      �?	             0@       ������������������������       �                     $@v      ������������������������       �r�q��?             @�      M       ^                 ��Y7@2�ߣ0��?Z            `a@      N       W                    �?П[;U��?9            �U@      O       R                    �?�X����?             F@       P       Q                 ��-@؇���X�?	             ,@       ������������������������       ����Q��?             @�       ������������������������       �                     "@      S       V                 03�1@���Q��?             >@      T       U                    �?      �?             4@       ������������������������       �      �?              @g      ������������������������       �      �?             (@�       ������������������������       �z�G�z�?             $@y       X       Y                    �?�K��&�?            �E@        ������������������������       ����Q��?             4@�       Z       ]                  �3@��+7��?             7@       [       \                    �?     ��?             0@       ������������������������       �z�G�z�?             $@        ������������������������       �r�q��?             @        ������������������������       �և���X�?             @        _       `                    �?4��?�?!             J@        ������������������������       ��q�q�?             @        a       b                    @��<b�ƥ?             G@        ������������������������       �      �?              @        ������������������������       �                     C@        �t�bh�h)h,K ��h.��R�(KKcKK��h\�B0       0|@     Pp@     `l@      M@      F@      ;@      A@      ;@       @      @      @@      4@      :@      @      @      �?      7@      @      "@      �?      ,@       @      @      0@      $@             �f@      ?@      d@      5@      L@      @     �A@      @      ;@      �?      *@              ,@      �?      @              @      �?       @       @      5@              Z@      2@      *@       @      @      @      @       @     �V@      $@      &@              T@      $@      7@      $@      ,@      "@       @       @      @      �?      "@      �?      l@     `i@      `@     �c@      D@      4@      B@      @      @      @      >@      @      &@      @      3@              @      ,@      @      @              $@     @V@     `a@      V@     �E@       @       @     �U@     �A@      S@     �A@      R@      9@      F@      5@      >@      1@      &@      ,@      3@      @      (@      �?      @      �?      @              @       @      ,@      @      <@      @      (@      @      @       @      @       @      0@              @      $@       @       @       @       @      $@              �?      X@             @T@      �?      .@              $@      �?      @     �W@      F@      H@     �C@      >@      ,@      (@       @      @       @      "@              2@      (@      $@      $@      @      �?      @      "@       @       @      2@      9@      (@       @      @      1@      @      *@       @       @      �?      @      @      @     �G@      @       @      @     �F@      �?      @      �?      C@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��nhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKihth)h,K ��h.��R�(KKi��h{�B@         R                  x#J@�"Y�\7�?�           @�@              	                    @<��Vi)�?~           ��@      �?                           �?\�Uo��?             C@ 0��  ������������������������       �                     &@�����                              @X�<ݚ�?             ;@      �?������������������������       �                     @                                   @      �?             4@      @������������������������       ��	j*D�?             *@      $@������������������������       �؇���X�?             @      �?
       +                 `f#@tTsy���?f           x�@      @       "                    �?��C��?�            �p@                               �?�@�Cc}h��?�             l@    `a@                          @@@P�� �?U            @`@    �A@                        �Y�@�$��y��?A            @X@      ,@                           �?�>4և��?             <@       ������������������������       �؇���X�?             ,@      @                        ��@d}h���?
             ,@       ������������������������       �                      @�      ������������������������       �      �?             @�      ������������������������       �p��%���?,            @Q@w      ������������������������       �                    �@@n                              ��y @Df/��?8            �W@                                �4@���y4F�?$            �L@       ������������������������       ��q�q�?             (@�                                �>@���V��?            �F@                                 ;@$�q-�?             :@       ������������������������       �                     $@      ������������������������       �      �?             0@                                �@@�d�����?             3@       ������������������������       ��q�q�?             @(      ������������������������       �$�q-�?             *@V              !                 ���"@�?�|�?            �B@      ������������������������       �                     :@3      ������������������������       ��C��2(�?             &@A      #       *                 @3�@      �?             D@       $       '                   �9@������?             >@        %       &                   �5@      �?
             0@       ������������������������       ����|���?             &@j       ������������������������       ����Q��?             @�       (       )                    �?؇���X�?
             ,@       ������������������������       �؇���X�?             @�       ������������������������       �؇���X�?             @�       ������������������������       ��z�G��?             $@$       ,       ?                    �?fܶ���?�            pr@       -       .                     �?,sI�v�?s            �f@        ������������������������       ��q�q�?"             H@-       /       0                 �&@�C��2(�?Q            �`@        ������������������������       �������?	             .@�       1       2                    �?|�űN�?H            @]@        ������������������������       ��<ݚ�?             "@�       3       >                    �?�X�<ݺ?A             [@       4       5                    �?�qM�R��?*            �P@        ������������������������       �����X�?             @�       6       ;                 039@��S�ۿ?%             N@      7       :                   �*@ �q�q�?             H@        8       9                   �=@ףp=
�?             4@       ������������������������       �                      @:      ������������������������       �r�q��?             (@;      ������������������������       �                     <@?      <       =                   @D@r�q��?             (@       ������������������������       �����X�?             @7      ������������������������       �                     @G       ������������������������       �                    �D@      @       A                   �0@84(���?K            �\@       ������������������������       ��8��8��?             (@�      B       G                     @ڲ�-���?D            �Y@      C       F                   �8@�O4R���?%            �J@        D       E                   �7@�C��2(�?	             &@      ������������������������       �                     @      ������������������������       �      �?             @-      ������������������������       �                     E@,      H       I                    �?�q�����?             I@       ������������������������       ��q�q�?             (@�       J       Q                 ���4@�\��N��?             C@       K       P                    �?X�Cc�?             <@      L       O                    @@�q�q�?             8@      M       N                    �?��S���?	             .@       ������������������������       ��z�G��?             $@�      ������������������������       �z�G�z�?             @�      ������������������������       ������H�?             "@�      ������������������������       �      �?             @�       ������������������������       �                     $@      S       \                    �?8����?I            �\@      T       U                   �3@�t����?)             Q@       ������������������������       �����X�?             @g      V       [                    �?\#r��?%            �N@        W       Z                     @d}h���?             <@       X       Y                    �?�z�G��?             4@        ������������������������       ��q�q�?             @�       ������������������������       �����X�?             ,@        ������������������������       �                      @        ������������������������       �                    �@@        ]       ^                 @3#O@�[�IJ�?             �G@        ������������������������       �                     @        _       h                    @X�Cc�?             E@       `       e                    �?�g�y��?             ?@       a       d                 03c@�E��ӭ�?             2@       b       c                 03�S@      �?             $@        ������������������������       �z�G�z�?             @        ������������������������       �z�G�z�?             @        ������������������������       �                      @        f       g                    <@�θ�?
             *@        ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                     &@        �t�bh�h)h,K ��h.��R�(KKiKK��h\�B�       �|@     `o@     �z@     `e@      .@      7@              &@      .@      (@              @      .@      @      "@      @      @      �?     �y@     �b@      k@     �G@     @i@      6@     @^@      "@      V@      "@      7@      @      (@       @      &@      @       @              @      @     @P@      @     �@@             @T@      *@     �F@      (@      @      @      C@      @      8@       @      $@              ,@       @      ,@      @       @      @      (@      �?      B@      �?      :@              $@      �?      .@      9@       @      6@      @      $@      @      @       @      @       @      (@      �?      @      �?      @      @      @     @h@     @Y@     �c@      6@      C@      $@      ^@      (@      &@      @     @[@       @      @       @     �Y@      @     �N@      @      @       @      L@      @      G@       @      2@       @       @              $@       @      <@              $@       @      @       @      @             �D@              B@     �S@      &@      �?      9@     �S@      �?      J@      �?      $@              @      �?      @              E@      8@      :@      @       @      4@      2@      $@      2@       @      0@      @       @      @      @      @      �?      �?       @       @       @      $@             �A@      T@       @      N@       @      @      @     �K@      @      6@      @      ,@       @      @      @      $@               @             �@@      ;@      4@              @      ;@      .@      0@      .@      *@      @      @      @      @      �?      �?      @       @              @      $@      @       @               @      &@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJXk�hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKkhth)h,K ��h.��R�(KKk��h{�B�         ,                     @��ے@R�?�           @�@                                   /@�r�����?�            Ps@      .@                           @�C��2(�?             6@        ������������������������       �����X�?             @      @������������������������       �        
             .@      @       !                  x#J@�!I���?�            �q@     @                           @�LQ�1	�?p             g@       @������������������������       �                     &@      �?	                        `f�:@NR�l���?i            �e@     6@
                          �*@     ��?N             `@      (@������������������������       � 1_#�?%            �M@     @Y@                           �?ꮃG��?)            @Q@     @                        ��D:@��s����?             E@     @                        03�9@h�����?             <@       @������������������������       �                     &@       @                           �?�IєX�?             1@    �S@������������������������       �                     "@Z      ������������������������       �      �?              @�      ������������������������       �      �?             ,@�                                 6@ 7���B�?             ;@       ������������������������       ��C��2(�?             &@n      ������������������������       �                     0@�                                  �?������?            �F@                                  �?:�&���?            �C@                                 �?��a�n`�?             ?@       ������������������������       �����X�?             @c                                �=@�q�q�?             8@                              ��yC@����X�?	             ,@      ������������������������       �և���X�?             @�      ������������������������       �                     @(      ������������������������       �ףp=
�?             $@V      ������������������������       �                      @J      ������������������������       �r�q��?             @3      "       +                    �?~�X��?A            �Y@       #       (                   �D@��V#�?            �E@       $       '                   �@@�q�����?             9@       %       &                    �?p�ݯ��?             3@       ������������������������       ��q�q�?             (@j       ������������������������       �����X�?             @�       ������������������������       �r�q��?             @�       )       *                 �UcV@�����H�?             2@       ������������������������       �      �?              @�       ������������������������       �                     $@$       ������������������������       �        #             N@       -       R                    �?h�*���?           0y@       .       /                    @�p�Ð�?�            Pq@        ������������������������       ����Q��?             $@]       0       7                    �?��c+��?�            �p@        1       6                    �?� ��1�?            �D@       2       3                 ���@��a�n`�?             ?@        ������������������������       �                     &@�       4       5                   @<@R���Q�?             4@       ������������������������       �8�Z$���?             *@�       ������������������������       �؇���X�?             @      ������������������������       �      �?             $@�       8       Q                 �T�I@�=|+g��?�            @l@      9       <                 ��@�n���?�             k@       :       ;                   �;@�q�q�?             (@       ������������������������       �և���X�?             @?      ������������������������       �                     @I      =       P                 ��y @�K��?�            �i@      >       O                    �?T�n��?X             b@       ?       B                   �:@�iyw	
�?T            �`@       @       A                   �2@�Ń��̧?             E@       ������������������������       �؇���X�?             @�      ������������������������       �                    �A@�      C       D                  s�@���}<S�?9             W@        ������������������������       �                     ,@8      E       J                   �?@��-�=��?1            �S@      F       I                   @@      �?             L@       G       H                 ��@���N8�?
             5@      ������������������������       �ףp=
�?             $@�      ������������������������       ����|���?             &@�       ������������������������       � >�֕�?            �A@�       K       L                 �?�@���7�?             6@       ������������������������       �        	             (@�      M       N                   �D@ףp=
�?	             $@      ������������������������       �                     @�      ������������������������       �      �?             @�      ������������������������       �z�G�z�?             $@�      ������������������������       �        +             N@�       ������������������������       �      �?             $@      S       X                    �?p<�w���?R            �_@       T       W                    �?�p ��?            �D@      U       V                 �&B@��a�n`�?             ?@      ������������������������       �؇���X�?             5@�       ������������������������       �                     $@y       ������������������������       ��z�G��?             $@}       Y       h                   �>@�ucQ?-�?7            @U@       Z       e                   �;@      �?,             Q@       [       ^                 pf� @��V#�?            �E@        \       ]                 �&B@��S���?             .@        ������������������������       �      �?              @        ������������������������       �և���X�?             @        _       d                    7@d}h���?             <@       `       c                    @��2(&�?             6@       a       b                    �?��S�ۿ?
             .@        ������������������������       ������H�?             "@        ������������������������       �                     @        ������������������������       �����X�?             @        ������������������������       �      �?             @        f       g                    �?H%u��?             9@        ������������������������       ����!pc�?             &@        ������������������������       �                     ,@        i       j                   @B@��.k���?             1@       ������������������������       ������H�?             "@        ������������������������       �      �?              @        �t�bh�h)h,K ��h.��R�(KKkKK��h\�B�       �|@     �o@     �b@     �c@       @      4@       @      @              .@     �b@     @a@      ^@      P@      &@             @[@      P@      S@      J@     �D@      2@     �A@      A@      A@       @      ;@      �?      &@              0@      �?      "@              @      �?      @      @      �?      :@      �?      $@              0@     �@@      (@      @@      @      8@      @      @       @      3@      @      $@      @      @      @      @              "@      �?       @              �?      @      =@     �R@      =@      ,@      *@      (@      (@      @      @      @      @       @      �?      @      0@       @      @       @      $@                      N@     @s@     �W@     `n@      A@      @      @     �m@      <@     �@@       @      <@      @      &@              1@      @      &@       @      @      �?      @      @     �i@      4@      i@      .@       @      @      @      @      @              h@      &@     �`@      &@     @_@      "@     �D@      �?      @      �?     �A@              U@       @      ,@             �Q@       @     �H@      @      0@      @      "@      �?      @      @     �@@       @      5@      �?      (@              "@      �?      @              @      �?       @       @      N@              @      @     @P@     �N@      @     �A@      @      <@      @      2@              $@      @      @     �M@      :@     �I@      1@      =@      ,@      @       @      @      @      @      @      6@      @      3@      @      ,@      �?       @      �?      @              @       @      @      @      6@      @       @      @      ,@               @      "@      �?       @      @      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ0��JhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKihth)h,K ��h.��R�(KKi��h{�B@         ,                     @�d��Pb�?�           @�@                                 x#J@~����m�?�            u@ be use                           �?\�����?�            �k@     G@                           (@z�c�@-�?a            �b@      (@������������������������       �                     @      :@                            �?:��o#@�?\            �a@      @                        `f�B@�̚��?'            �N@     @                           B@֭��F?�?            �G@        	                           =@      �?             2@     (@
                        �ܵ<@�q�q�?
             (@      @������������������������       �z�G�z�?             @      N@������������������������       �և���X�?             @      <@������������������������       ��q�q�?             @      @                          �G@8^s]e�?             =@      4@                        03k:@r�q��?             (@        ������������������������       �؇���X�?             @      �?������������������������       �z�G�z�?             @Z                                 <@j���� �?	             1@      ������������������������       �      �?              @�      ������������������������       �X�<ݚ�?             "@w      ������������������������       �                     ,@n                                 �?ףp=
�?5             T@                                �;@Ԫ2��?'            �L@       ������������������������       ����N8�?             5@�      ������������������������       �tk~X��?             B@�      ������������������������       �                     7@c                                 6@�k~X��?(             R@                                  �?г�wY;�?             A@      ������������������������       �                     7@�      ������������������������       ��C��2(�?             &@(      ������������������������       �                     C@V              +                    �?��Sݭg�?E            @]@       !       $                    �?j���� �?            �I@       "       #                    �?�G��l��?
             5@      ������������������������       ��C��2(�?             &@�       ������������������������       �ףp=
�?             $@�       %       *                    �?�q�q�?             >@       &       '                 ��,P@�q�q�?             8@        ������������������������       ����Q��?             @�       (       )                   �D@�KM�]�?
             3@       ������������������������       �                     (@�       ������������������������       �����X�?             @�       ������������������������       �r�q��?             @$       ������������������������       �        )            �P@       -       2                    @b����o�?�            pw@        .       1                 03�9@�5��?             ;@       /       0                    �?      �?
             0@        ������������������������       �r�q��?             @�       ������������������������       �                     $@A       ������������������������       ��C��2(�?             &@�       3       X                 ��.@��&y�X�?�            �u@       4       U                    �?��{H�?�            Pp@       5       P                    �?�֪u�_�?�            �m@       6       K                   @@@,���$�?}            @h@      7       J                   �?@ghډC�?_            �b@       8       ?                   �;@,�d�vK�?Z            �a@       9       >                   �8@h��@D��?,            �Q@      :       =                   �4@�X�<ݺ?&             K@      ;       <                 pf� @�����H�?             ;@      ������������������������       �     ��?             0@I      ������������������������       �                     &@7      ������������������������       �                     ;@G       ������������������������       �������?             1@      @       I                   �<@����Q8�?.            �Q@      A       H                 ��) @Hn�.P��?(             O@      B       G                 �?$@ 7���B�?!             K@      C       F                    �?@4և���?             <@       D       E                 ���@���7�?             6@       ������������������������       �ףp=
�?             $@      ������������������������       �                     (@-      ������������������������       �r�q��?             @,      ������������������������       �                     :@�      ������������������������       �      �?              @�       ������������������������       ������H�?             "@�       ������������������������       �      �?              @v      L       M                   �E@`���i��?             F@      ������������������������       �                     =@�      N       O                 ��Y@��S�ۿ?             .@      ������������������������       �                     @�      ������������������������       �      �?              @�      Q       T                 ���@X�Cc�?             E@        R       S                   �3@      �?             0@       ������������������������       �r�q��?             @-      ������������������������       �                     $@%      ������������������������       ���
ц��?             :@g      V       W                    �?`2U0*��?             9@       ������������������������       �                     5@y       ������������������������       �      �?             @}       Y       d                 03�7@8^s]e�?:            �U@        Z       c                   @@@z�J��?            �G@       [       `                    �?b�2�tk�?             B@       \       _                    �?�㙢�c�?             7@       ]       ^                    ;@�t����?             1@        ������������������������       �      �?             @        ������������������������       �$�q-�?             *@        ������������������������       ��q�q�?             @        a       b                    �?�θ�?
             *@        ������������������������       �؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �"pc�
�?             &@        e       h                    �?ףp=
�?             D@        f       g                 0�H@���|���?             &@        ������������������������       �                     @        ������������������������       �z�G�z�?             @        ������������������������       �                     =@        �t�b��     h�h)h,K ��h.��R�(KKiKK��h\�B�       @{@     @q@     @b@     �g@      ]@      Z@     �\@     �@@              @     �\@      :@     �E@      2@      =@      2@      "@      "@      @      @      @      �?      @      @       @      @      4@      "@      $@       @      @      �?      @      �?      $@      @      @      @      @      @      ,@              R@       @     �H@       @      4@      �?      =@      @      7@              �?     �Q@      �?     �@@              7@      �?      $@              C@      >@     �U@      >@      5@      $@      &@      �?      $@      "@      �?      4@      $@      3@      @       @      @      1@       @      (@              @       @      �?      @             �P@      r@     @U@      &@      0@      �?      .@      �?      @              $@      $@      �?     pq@     @Q@     `k@      E@     `h@     �D@     �f@      ,@      a@      *@     ``@      &@      P@      @     �I@      @      8@      @      *@      @      &@              ;@              *@      @     �P@      @     �M@      @      J@       @      :@       @      5@      �?      "@      �?      (@              @      �?      :@              @      �?       @      �?      @       @     �E@      �?      =@              ,@      �?      @              @      �?      .@      ;@      �?      .@      �?      @              $@      ,@      (@      8@      �?      5@              @      �?      N@      ;@      8@      7@      6@      ,@      3@      @      .@       @      @      �?      (@      �?      @       @      @      $@      �?      @       @      @       @      "@      B@      @      @      @      @              �?      @      =@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJڡWhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKghth)h,K ��h.��R�(KKg��h{�B�         X                  x#J@�1�uџ�?�           @�@              =                    �?�z��U�?t           p�@     2@                           @v^|�_�?           �z@      �?                           �?���!pc�?             &@        ������������������������       �                     @      @������������������������       �      �?             @      �?       ,                   �A@j:?���?           �y@    �@@       +                    @r�q��?�            �s@    �U@	       
                    ,@���I��?�            �r@      �?������������������������       �r�q��?             @       @       &                   �?@ZՏ�m|�?�            `r@    �P@       %                    �?R��q�?�             p@     @       $                    �?4?,R��?�            �o@     E@       !                    �?���!�=�?�            �n@     &@                           �?�
���?�             k@      @                           ;@д>��C�?             =@      @������������������������       ����Q��?             @Z                              ��%@      �?             8@      ������������������������       �      �?             0@�      ������������������������       �      �?              @w                                 @@ l{wY|�?y            �g@                                   @H�V�e��?'             Q@       ������������������������       �                     &@�                              ��@P̏����?!            �L@                                 7@:�&���?            �C@       ������������������������       �                     @c                              ���@�'�`d�?            �@@       ������������������������       �X�<ݚ�?             "@      ������������������������       �      �?             8@�                                �:@b�2�tk�?             2@       ������������������������       ��q�q�?             "@V      ������������������������       �X�<ݚ�?             "@J      ������������������������       �2Tv���?R             ^@3      "       #                 ��l#@ܷ��?��?             =@       ������������������������       ��q�q�?             "@�       ������������������������       �                     4@�       ������������������������       �                     @v       ������������������������       �      �?             @j       '       (                     @�E��ӭ�?             B@        ������������������������       ��ՙ/�?             5@�       )       *                 @3�@�r����?             .@       ������������������������       �      �?              @�       ������������������������       �                     @$       ������������������������       �                     2@       -       6                 ��$:@DE�SA_�?;            @X@       .       5                    �?F��}��?)            @R@       /       0                     @����?%            @P@        ������������������������       �ܷ��?��?             =@�       1       2                    �?������?             B@        ������������������������       �                     @�       3       4                 pff@      �?             @@       ������������������������       �        
             1@�       ������������������������       ���S�ۿ?             .@�       ������������������������       �                      @      7       <                   �L@r�q��?             8@       8       9                 `f&;@      �?             0@       ������������������������       �      �?             @:      :       ;                    G@�8��8��?	             (@      ������������������������       �                     @?      ������������������������       �z�G�z�?             @I      ������������������������       �                      @7      >       A                     @�=���D�?f            �d@        ?       @                    �?p���?             I@       ������������������������       �ףp=
�?             $@!      ������������������������       �                     D@�      B       S                    �?`3�a���?G            �\@      C       R                 ��*4@      �?7             V@       D       Q                    .@=&C��?3            �T@      E       P                    �?<��¤�?+             Q@      F       I                    �?��۾%d�?%             M@       G       H                 ��@�X����?             6@      ������������������������       ��r����?             .@�      ������������������������       �����X�?             @�       J       O                 ��i#@      �?             B@       K       N                   �;@*;L]n�?             >@      L       M                 �&B@������?	             .@      ������������������������       �      �?              @�      ������������������������       �؇���X�?             @�      ������������������������       ����Q��?             .@�      ������������������������       �r�q��?             @�      ������������������������       �z�G�z�?             $@�       ������������������������       ��r����?             .@      ������������������������       �z�G�z�?             @-      T       U                 `v�6@�θ�?             :@       ������������������������       �����X�?             @g      V       W                 ��T?@�}�+r��?             3@        ������������������������       �                     (@y       ������������������������       �؇���X�?             @}       Y       d                    �?ҐϿ<��?O            �^@        Z       _                 Ј�U@��U/��?&            �L@       [       \                   �;@�n`���?             ?@        ������������������������       �      �?              @        ]       ^                    �?���}<S�?             7@        ������������������������       ��q�q�?             @        ������������������������       �                     1@        `       c                    �?
j*D>�?             :@       a       b                  ��^@      �?
             0@       ������������������������       ��q�q�?             "@        ������������������������       �؇���X�?             @        ������������������������       ��z�G��?             $@        e       f                    �?��ɉ�?)            @P@       ������������������������       �        "            �L@        ������������������������       �      �?              @        �t�bh�h)h,K ��h.��R�(KKgKK��h\�Bp       P|@     0p@     �y@     `f@     Pv@     @Q@      @       @              @      @      �?      v@     �N@     �p@     �J@     �n@     �J@      �?      @     �n@      H@     �k@      C@      k@     �A@     `j@     �A@      g@      @@      8@      @      @       @      5@      @      .@      �?      @       @      d@      ;@      K@      ,@      &@             �E@      ,@      @@      @      @              :@      @      @      @      5@      @      &@      @      @      @      @      @     �Z@      *@      :@      @      @      @      4@              @              @      @      :@      $@      *@       @      *@       @      @       @      @              2@             @V@       @     @Q@      @     �N@      @      :@      @     �A@      �?      @              ?@      �?      1@              ,@      �?       @              4@      @      (@      @      �?      @      &@      �?      @              @      �?       @              K@     �[@      �?     �H@      �?      "@              D@     �J@     �N@     �@@     �K@      =@      K@      ;@     �D@      9@     �@@      @      .@       @      *@      @       @      2@      2@      *@      1@      @      &@      @      @      �?      @      "@      @      @      �?       @       @       @      *@      @      �?      4@      @       @      @      2@      �?      (@              @      �?      E@      T@      D@      1@      9@      @      @      @      5@       @      @       @      1@              .@      &@      (@      @      @      @      @      �?      @      @       @     �O@             �L@       @      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ:d�hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKghth)h,K ��h.��R�(KKg��h{�B�         @                    �?���x�W�?�           @�@              '                 039@���J��?           �{@     @                            �?����
R�?�            �s@     ,@       	                    �?dP-���?�            �q@      @                          �=@r�q��?             >@      @                        ��%@��<b���?             7@     ,@������������������������       �����X�?             ,@      @������������������������       ������H�?             "@      @������������������������       �                     @        
                           �?�����?�            �o@      @                          �0@��Au5a�?�            �k@        ������������������������       �      �?              @      @                          �<@����Q8�?�            �j@                               �?$@��.N"Ҭ?V            @a@      @                         s�@$�q-�?            �C@     �?                           �? 7���B�?             ;@      "@������������������������       �                     @Z                              @33@P���Q�?             4@       ������������������������       �ףp=
�?             $@�      ������������������������       �                     $@w                              ��@r�q��?	             (@      ������������������������       �r�q��?             @�      ������������������������       �r�q��?             @�                              ���$@`�LVXz�?<            �X@      ������������������������       �        )            @Q@�                                �(@(;L]n�?             >@       ������������������������       �؇���X�?             @      ������������������������       �                     7@                                  @H0sE�d�?1            �R@       ������������������������       ��r����?	             .@(      ������������������������       �ףp=
�?(             N@V      ������������������������       ��חF�P�?             ?@J      !       $                 �y�/@*O���?             B@       "       #                    ;@��.k���?
             1@      ������������������������       �      �?             (@�       ������������������������       �                     @�       %       &                    #@���y4F�?             3@        ������������������������       �z�G�z�?             @j       ������������������������       �                     ,@�       (       +                    �?b �y��?S            �_@        )       *                    �?�g�y��?             ?@       ������������������������       �X�<ݚ�?             2@�       ������������������������       ���
ц��?             *@$       ,       1                   �>@�q�q�?A             X@        -       0                     �?`՟�G��?             ?@       .       /                   �A@j���� �?             1@        ������������������������       �      �?             @]       ������������������������       ��	j*D�?             *@�       ������������������������       �����X�?
             ,@A       2       3                    @&����?+            @P@        ������������������������       ����Q��?             @�       4       7                  x#J@���*�?'             N@        5       6                    $@ ��WV�?             :@        ������������������������       �؇���X�?             @      ������������������������       �                     3@�       8       ;                 �!�N@�t����?             A@       9       :                      @���Q��?             $@       ������������������������       ��q�q�?             @;      ������������������������       �                     @?      <       ?                    @r�q��?             8@      =       >                    �?      �?
             0@      ������������������������       ��z�G��?             $@G       ������������������������       �r�q��?             @      ������������������������       �                      @!      A       L                     @���Őm�?�            �p@      B       K                 03[=@��.N"Ҭ?U            @a@       C       D                     �?����Q8�?(            �Q@        ������������������������       �և���X�?             @8      E       J                   �;@     ��?$             P@       F       G                   �3@ �q�q�?             8@       ������������������������       �                     *@,      H       I                    �?�C��2(�?	             &@       ������������������������       �                     @�       ������������������������       �z�G�z�?             @�       ������������������������       �                     D@v      ������������������������       �        -            �P@�      M       \                    �?v ��?P             `@      N       Q                 ���@b1<+�C�?1            @R@       O       P                 P�@     ��?             0@      ������������������������       ����!pc�?             &@�      ������������������������       �                     @�       R       W                    �?T�7�s��?&            �L@      S       V                 pF @      �?             C@      T       U                   �6@���|���?             6@       ������������������������       �؇���X�?             @g      ������������������������       ���S���?
             .@�       ������������������������       �     ��?             0@y       X       Y                    �?�����?             3@        ������������������������       �z�G�z�?             @�       Z       [                 ��80@X�Cc�?             ,@        ������������������������       �և���X�?             @        ������������������������       �؇���X�?             @        ]       d                    �?���X�?             L@       ^       _                    �?�q�q�?             B@        ������������������������       ����Q��?             $@        `       c                   �>@�θ�?             :@       a       b                    �?P���Q�?	             4@       ������������������������       �؇���X�?             @        ������������������������       �                     *@        ������������������������       �r�q��?             @        e       f                    @R���Q�?             4@        ������������������������       �      �?             @        ������������������������       �        	             ,@        �t�bh�h)h,K ��h.��R�(KKgKK��h\�Bp       P{@     0q@     �v@     @T@     �q@     �B@      p@      8@      9@      @      2@      @      $@      @       @      �?      @              m@      3@     �i@      ,@      @       @      i@      (@     �`@      @      B@      @      :@      �?      @              3@      �?      "@      �?      $@              $@       @      @      �?      @      �?     �X@      �?     @Q@              =@      �?      @      �?      7@             �P@       @      *@       @      K@      @      :@      @      7@      *@       @      "@      @      "@      @              .@      @      �?      @      ,@             �T@      F@      .@      0@       @      $@      @      @      Q@      <@      1@      ,@      @      $@      @      �?      @      "@      $@      @     �I@      ,@       @      @     �H@      &@      9@      �?      @      �?      3@              8@      $@      @      @      @       @              @      4@      @      (@      @      @      @      @      �?       @             @R@     @h@      @     �`@      @     �P@      @      @      �?     �O@      �?      7@              *@      �?      $@              @      �?      @              D@             �P@     @Q@      N@      <@     �F@      @      *@      @       @              @      9@      @@      3@      3@       @      ,@      �?      @      @       @      &@      @      @      *@      �?      @      @      "@      @      @      �?      @     �D@      .@      8@      (@      @      @      4@      @      3@      �?      @      �?      *@              �?      @      1@      @      @      @      ,@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�I]fhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK
hsKUhth)h,K ��h.��R�(KKU��h{�B@         6                    �?������?�           @�@                                  @X�'�f��?            }@      �?                            @ҳ�wY;�?             A@        ������������������������       �                     &@                                ���8@
;&����?             7@        ������������������������       �                     $@      �?������������������������       �$�q-�?             *@                                  �5@���tT��?           �z@      @	                           �?�>����?/            @T@       
                          �2@����˵�?!            �M@      F@������������������������       �                     7@      <@                          �3@�8��8��?             B@      "@������������������������       �d}h���?             ,@      &@������������������������       �                     6@      $@                            @��2(&�?             6@      @������������������������       �      �?             @                                ��A>@�X�<ݺ?
             2@       ������������������������       �      �?              @�      ������������������������       �                     $@�             !                     �?\�&�s��?�            �u@                                 @B@>��C��?2            �U@                               Ј�Q@�G�z�?             D@      ������������������������       �d}h���?             <@�      ������������������������       ��q�q�?             (@�                                �E@*
;&���?             G@                              ��>@�GN�z�?             6@                                 J@�r����?
             .@       ������������������������       �����X�?             @      ������������������������       �                      @�      ������������������������       �և���X�?             @(                                 @G@�8��8��?             8@       ������������������������       �                     &@J      ������������������������       �8�Z$���?             *@3      "       5                 0��G@�~�H��?�            pp@      #       *                 �Y�@$%j����?�            �o@        $       %                   �;@z�G�z�?            �A@        ������������������������       �      �?              @v       &       )                    �? 7���B�?             ;@        '       (                 ���@�C��2(�?	             &@       ������������������������       �                     @�       ������������������������       �      �?             @�       ������������������������       �        
             0@�       +       4                    �?��<nd�?�            @k@       ,       -                 @3�@TxH���?�            �j@        ������������������������       ������H�?4            �V@       .       1                     @�&/�E�?U             _@        /       0                   �;@�*/�8V�?#            �G@        ������������������������       �        	             *@�       ������������������������       ���hJ,�?             A@A       2       3                    �?�g<a�?2            @S@        ������������������������       �r�q��?             (@�       ������������������������       �        +            @P@�       ������������������������       �      �?             @�       ������������������������       ����Q��?             $@      7       >                     @�y��A�?�             o@       8       9                    @�J�T�?X            �a@       ������������������������       �      �?              @:      :       ;                    �? 
�V�?T            �`@      ������������������������       �        E            �[@?      <       =                 ���`@ �q�q�?             8@      ������������������������       �                     0@7      ������������������������       �      �?              @G       ?       T                 `v�6@�����?@            �Z@      @       G                    �?ܐ҆��?6            @W@       A       D                 P��+@�����?             C@      B       C                  s�@R���Q�?             4@       ������������������������       ����Q��?             @8       ������������������������       �        	             .@8      E       F                    �?      �?             2@       ������������������������       �      �?              @-      ������������������������       ����Q��?             $@,      H       M                   �6@N{�T6�?!            �K@       I       L                    �?�q�q�?             8@       J       K                   �4@����X�?             ,@        ������������������������       ����Q��?             @v      ������������������������       ��<ݚ�?             "@�      ������������������������       �ףp=
�?             $@�      N       S                 ��Y.@�g�y��?             ?@      O       P                   �;@�E��ӭ�?             2@       ������������������������       �և���X�?             @�      Q       R                   #@�C��2(�?             &@        ������������������������       �                     @      ������������������������       �z�G�z�?             @-      ������������������������       �8�Z$���?             *@%      ������������������������       �        
             *@g      �t�bh�h)h,K ��h.��R�(KKUKK��h\�BP        |@     `p@     0x@     @S@      (@      6@              &@      (@      &@              $@      (@      �?     pw@     �K@     �R@      @      L@      @      7@             �@@      @      &@      @      6@              3@      @       @       @      1@      �?      @      �?      $@             �r@     �H@     �P@      4@      ;@      *@      6@      @      @      @     �C@      @      1@      @      *@       @      @       @       @              @      @      6@       @      &@              &@       @     @m@      =@     �l@      9@      <@      @       @      @      :@      �?      $@      �?      @              @      �?      0@              i@      2@     �h@      1@      T@      $@     @]@      @      E@      @      *@              =@      @     �R@       @      $@       @     @P@              @      �?      @      @     �O@      g@      @     @a@      @      @      �?     �`@             �[@      �?      7@              0@      �?      @     �M@     �G@      G@     �G@      (@      :@      @      1@      @       @              .@      "@      "@      @      @      @      @      A@      5@      3@      @      $@      @      @       @      @       @      "@      �?      .@      0@      *@      @      @      @      $@      �?      @              @      �?       @      &@      *@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�޵#hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKshth)h,K ��h.��R�(KKs��h{�B�         ^                 `f~I@~�Я��?�           @�@                                  !@��}y.��?e           ȁ@     �K@                           @�I� �?             G@     (@������������������������       �                     <@       @                        ��T?@r�q��?             2@    �H@������������������������       �                     (@      @������������������������       �      �?             @       @       ?                    �? �&4��?H           X�@       	       8                 ��$:@�LQ�1	�?�             w@     @
       7                 ��Y7@�4�?�            ps@                                 �0@P�I;l�?�            �q@      1@������������������������       �      �?              @               6                 0#�2@䦳	�R�?�            0q@              5                 `��+@(�=�]�?�            �p@    @a@                            @����2�?�             n@      7@                          �@@>a�����?            �I@    �G@                           ;@�C��2(�?            �@@ �ex�7                          �'@      �?             0@ ���H�������������������������       �ףp=
�?             $@/����L������������������������       �                     @��̔׾�                        `fF)@�t����?             1@6m��R\������������������������       �                     (@�33���C�������������������������       ����Q��?             @n��Y���                        ��Y)@�E��ӭ�?
             2@ v-b%��������������������������       �      �?              @���W�gd������������������������       ��z�G��?             $@�esU��J�                          �@�����H�?|            �g@ �\��i��������������������������       ����Q��?             @^�pu!�Q       0                 @3�@�_�����?x             g@��:^��       #                    �?��Ͻ��?W            @a@ ��GC                            �?������?            �D@ �"#h"�������������������������       ��IєX�?             1@�T�΀y��!       "                   �<@ �q�q�?             8@      ������������������������       �                     3@A      ������������������������       �z�G�z�?             @�       $       -                   @@@B�1V���?<            @X@       %       ,                 �?�@��G���?-            �R@       &       '                   �:@8�Z$���?(            @P@       ������������������������       �P���Q�?             D@�       (       +                   �@`�Q��?             9@       )       *                 ���@և���X�?	             ,@       ������������������������       �����X�?             @�       ������������������������       �؇���X�?             @$       ������������������������       �                     &@       ������������������������       �X�<ݚ�?             "@       .       /                  sW@�nkK�?             7@       ������������������������       �        
             0@]       ������������������������       �؇���X�?             @�       1       4                 0S�"@�nkK�?!             G@       2       3                    ?@�(\����?             D@       ������������������������       �                     :@�       ������������������������       �@4և���?
             ,@�       ������������������������       �r�q��?             @�       ������������������������       �XB���?             =@      ������������������������       ��q�q�?             @�       ������������������������       �                     <@`      9       >                 �D B@���y4F�?!            �L@      :       =                   `G@4�B��?            �B@      ;       <                   @C@ �o_��?             9@      ������������������������       �b�2�tk�?             2@I      ������������������������       �                     @7      ������������������������       ��q�q�?             (@G       ������������������������       �        
             4@      @       G                     @�y��<��?c            `c@       A       F                    6@X�EQ]N�?            �E@       B       C                 `f�)@z�G�z�?             9@       ������������������������       �                     $@8       D       E                   �<@�q�q�?
             .@       ������������������������       �����X�?             @      ������������������������       �                      @-      ������������������������       �                     2@,      H       [                    �?~h����?E             \@      I       J                 �&�@tv?z���?6            �V@        ������������������������       �                     @�       K       X                    .@Zz�����?2            @U@      L       Q                 pF @V{q֛w�?$             O@      M       N                   �9@և���X�?            �A@       ������������������������       �և���X�?	             ,@�      O       P                    �?�q�q�?
             5@      ������������������������       �      �?             (@�      ������������������������       ������H�?             "@�       R       S                 @33"@������?             ;@       ������������������������       �                     $@-      T       U                   �3@j���� �?             1@       ������������������������       ��q�q�?             @g      V       W                    =@���!pc�?	             &@        ������������������������       �r�q��?             @y       ������������������������       ����Q��?             @}       Y       Z                 ���6@�LQ�1	�?             7@       ������������������������       �@�0�!��?
             1@        ������������������������       �r�q��?             @        \       ]                 ��*4@�X����?             6@        ������������������������       ��z�G��?             $@        ������������������������       �        	             (@        _       l                    �?OX���?W            �a@        `       c                 03�M@�ʻ����?*             Q@        a       b                 �TL@������?             .@       ������������������������       �      �?              @        ������������������������       �؇���X�?             @        d       i                    �?H(���o�?            �J@        e       f                   �?@
;&����?             7@        ������������������������       ��q�q�?             (@        g       h                    �?���!pc�?             &@        ������������������������       �      �?             @        ������������������������       �؇���X�?             @        j       k                  D0T@�������?             >@       ������������������������       �        
             3@        ������������������������       ����|���?             &@        m       r                   �<@���Lͩ�?-            �R@        n       o                    �?z�G�z�?            �A@        ������������������������       �                     "@        p       q                 ���S@R�}e�.�?             :@        ������������������������       �      �?             $@        ������������������������       �      �?             0@        ������������������������       �                     D@        �t�bh�h)h,K ��h.��R�(KKsKK��h\�B0       �{@     �p@     �x@     `e@      .@      ?@              <@      .@      @      (@              @      @     �w@     �a@      t@      H@     0q@      B@     �n@      B@      @      @     `n@      @@     �m@      >@     `j@      =@     �E@       @      >@      @      .@      �?      "@      �?      @              .@       @      (@              @       @      *@      @      @       @      @      @      e@      5@      @       @     �d@      3@     @^@      1@     �C@       @      0@      �?      7@      �?      3@              @      �?     �T@      .@      N@      ,@     �K@      $@      C@       @      1@       @      @       @      @       @      �?      @      &@              @      @      6@      �?      0@              @      �?      F@       @     �C@      �?      :@              *@      �?      @      �?      <@      �?      @       @      <@             �F@      (@      9@      (@      2@      @      &@      @      @              @      @      4@             �O@      W@      @      C@      @      4@              $@      @      $@      @       @               @              2@      M@      K@     �E@     �G@              @     �E@      E@     �A@      ;@      .@      4@       @      @      @      ,@      @      @      �?       @      4@      @      $@              $@      @       @      @       @      @      @      �?      @       @       @      .@      @      ,@      @      �?      .@      @      @      @      (@             �F@     �X@      C@      >@      @      &@      @      @      �?      @      A@      3@      &@      (@       @      @      @       @       @       @      �?      @      7@      @      3@              @      @      @      Q@      @      <@              "@      @      3@      @      @       @      ,@              D@�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�G�hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKohth)h,K ��h.��R�(KKo��h{�B�         (                     @z����?�           @�@                                   �?B�F<��?�             s@                                  �?d���r��?�            �j@     1@       	                    �?������?U            @a@                                 �d@@�q�q�?             8@                                 �<@��S�ۿ?             .@      @������������������������       �      �?              @       @������������������������       �                     @      �?������������������������       ��q�q�?             "@      .@
                            �?�S����?G            �\@       @                        `f�;@�������?"             N@                                   G@8�A�0��?             6@     �?������������������������       ��q�q�?             (@      �?������������������������       �z�G�z�?             $@                                  �G@�?�'�@�?             C@     @                          �@@�>����?             ;@     W@                          �<@r�q��?	             (@       ������������������������       �z�G�z�?             @�      ������������������������       �؇���X�?             @�      ������������������������       �                     .@w      ������������������������       ����!pc�?             &@n      ������������������������       ��>����?%             K@�                                �6@�}�+r��?3             S@                                 �;@�J�4�?             9@       ������������������������       �����X�?             ,@�      ������������������������       �        	             &@c      ������������������������       �        #            �I@             !                   �8@$�ݏ^��?5            �V@                                 �2@ �#�Ѵ�?            �E@      ������������������������       �                     :@(                                  7@�t����?	             1@       ������������������������       ��q�q�?             @J      ������������������������       �                     &@3      "       %                    �?�[�IJ�?            �G@       #       $                    �? ��WV�?             :@        ������������������������       �                     ,@�       ������������������������       ��8��8��?             (@v       &       '                 pf�\@�����?             5@       ������������������������       �        
             ,@�       ������������������������       �����X�?             @�       )       4                    �?B(����?           �y@        *       3                 ���.@Ɣ��Hr�?'            �M@       +       ,                    0@�7����?            �G@        ������������������������       �����X�?             @       -       2                 �� @z�G�z�?             D@       .       1                    ?@r֛w���?             ?@       /       0                   �:@�q�q�?             8@        ������������������������       �����X�?             @�       ������������������������       �ҳ�wY;�?
             1@A       ������������������������       �                     @�       ������������������������       �                     "@�       ������������������������       �r�q��?             (@�       5       ^                    �?V�:וd�?�            �u@       6       9                    @�'F����?�            �o@       7       8                    �?     ��?             0@        ������������������������       �և���X�?             @`      ������������������������       �X�<ݚ�?             "@:      :       ]                    �?$�� ���?�            �m@      ;       \                 0�H@؇���X�?�            �l@      <       W                 ��i @`�t�D7�?�            �k@      =       N                 �?�@R�(CW�?d            �d@      >       M                   @@@�?�P�a�?G             ^@       ?       @                    �?8��8���?8             X@       ������������������������       �`Jj��?             ?@!      A       F                   �7@�����D�?(            @P@       B       E                 ��L@`2U0*��?             9@      C       D                   �5@$�q-�?	             *@        ������������������������       �r�q��?             @8      ������������������������       �                     @      ������������������������       �                     (@-      G       L                   �@��Q���?             D@      H       I                 ���@� �	��?             9@       ������������������������       �z�G�z�?             @�       J       K                   �:@��Q��?             4@        ������������������������       �r�q��?             @v      ������������������������       �և���X�?             ,@�      ������������������������       �        
             .@�      ������������������������       �                     8@�      O       T                    ?@���!pc�?             F@      P       Q                   �5@8�Z$���?             :@       ������������������������       �և���X�?             @�       R       S                    ;@�}�+r��?             3@       ������������������������       �                     @-      ������������������������       ��8��8��?	             (@%      U       V                 @3�@X�<ݚ�?
             2@       ������������������������       �      �?              @�       ������������������������       �z�G�z�?             $@y       X       Y                    )@XB���?*             M@        ������������������������       �z�G�z�?             @�       Z       [                    �?�O4R���?&            �J@       ������������������������       �                     ?@        ������������������������       ����7�?             6@        ������������������������       �X�<ݚ�?             "@        ������������������������       �                     @        _       `                  s�@���̅��?:            �W@        ������������������������       �                     $@        a       d                    �?���Q��?5            @U@        b       c                 03�'@��Q��?             4@       ������������������������       ���
ц��?             *@        ������������������������       �                     @        e       j                    �?@i��M��?*            @P@       f       i                    �?      �?             D@       g       h                   �9@�z�G��?             >@       ������������������������       �r�q��?	             2@        ������������������������       �      �?             (@        ������������������������       ����Q��?             $@        k       l                    �?�+e�X�?             9@        ������������������������       �և���X�?             @        m       n                    @r�q��?             2@       ������������������������       �                     "@        ������������������������       ��q�q�?             "@        �t�bh�h)h,K ��h.��R�(KKoKK��h\�B�       �{@     �p@     @b@     �c@     @]@     @X@     @\@      9@      1@      @      ,@      �?      @      �?      @              @      @      X@      2@      G@      ,@      *@      "@      @      @       @       @     �@@      @      9@       @      $@       @      @      �?      @      �?      .@               @      @      I@      @      @      R@      @      5@      @      $@              &@             �I@      =@     �N@       @     �D@              :@       @      .@       @      @              &@      ;@      4@      9@      �?      ,@              &@      �?       @      3@              ,@       @      @     �r@     �Z@      B@      7@      A@      *@       @      @      @@       @      7@       @      0@       @      @       @      &@      @      @              "@               @      $@     �p@      U@     �j@      D@      "@      @      @      @      @      @     �i@     �@@     �h@     �@@     @h@      <@     @a@      :@     �Z@      ,@     �T@      ,@      =@       @     �J@      (@      8@      �?      (@      �?      @      �?      @              (@              =@      &@      ,@      &@      �?      @      *@      @      @      �?       @      @      .@              8@              @@      (@      6@      @      @      @      2@      �?      @              &@      �?      $@       @       @      @       @       @      L@       @      @      �?      J@      �?      ?@              5@      �?      @      @      @             �I@      F@              $@     �I@      A@      @      *@      @      @              @      F@      5@      9@      .@      5@      "@      .@      @      @      @      @      @      3@      @      @      @      .@      @      "@              @      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ���JhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsK]hth)h,K ��h.��R�(KK]��h{�B@         *                     @�VM�?�           @�@                                   �?T �����?�             s@                               ��D:@f�B���?u            �i@      �?                           1@�ܸb���?4             W@ -}��  ������������������������       �z�G�z�?             @                                    �?X��%�?0            �U@      5@������������������������       �                      @     �N@������������������������       �86��Z�?,            �S@      @	                        ���X@����X�?A             \@       
                          �;@�~�����?8            �X@      @                        h"P@և���X�?
             ,@     @������������������������       ��z�G��?             $@       @������������������������       �      �?             @      $@                        ���S@���mC�?.            @U@     @                          �L@�<ݚ�?(             R@     <@                        ��";@r֛w���?!             O@       @������������������������       �z�G�z�?             @Z                                �<@���y4F�?            �L@                               `f�B@      �?
             0@      ������������������������       ��eP*L��?             &@w      ������������������������       �                     @n                                 �?�p ��?            �D@                                 �?      �?             @@       ������������������������       ��q�q�?             (@�      ������������������������       �        
             4@�      ������������������������       ��<ݚ�?             "@c      ������������������������       �                     $@      ������������������������       ���
ц��?             *@                                 �?$�q-�?	             *@       ������������������������       �                     @(      ������������������������       �؇���X�?             @V              !                    @г�wY;�?A            �Y@       ������������������������       �z�G�z�?             @3      "       '                   �H@`�E���?=            @X@      #       &                   �;@@�z�G�?3             T@        $       %                    6@�nkK�?             7@        ������������������������       �z�G�z�?             @v       ������������������������       �                     2@j       ������������������������       �        #            �L@�       (       )                     �?�IєX�?
             1@       ������������������������       �      �?              @�       ������������������������       �                     "@�       +       V                 ��Y7@���n�?�            `y@       ,       ;                    �?�c�x��?�            @u@        -       4                    �?���B��?@             [@       .       1                    ;@<���D�?(            �P@        /       0                   �4@����X�?
             ,@        ������������������������       ��q�q�?             @�       ������������������������       �      �?              @A       2       3                   �<@$�q-�?             J@       ������������������������       �                    �@@�       ������������������������       ����y4F�?             3@�       5       6                   �2@r�q��?             E@        ������������������������       �                     @      7       :                    �?tk~X��?             B@       8       9                 �&B@д>��C�?             =@      ������������������������       ��q�q�?	             .@:      ������������������������       �                     ,@;      ������������������������       �����X�?             @?      <       G                   �;@�EC�?�             m@       =       F                   @1@�(�Tw��?G            @]@      >       E                   �:@>�Q��?@             Z@       ?       @                    '@ʂy��?<            @X@       ������������������������       �      �?              @!      A       B                    �?��~l�?7            @V@      ������������������������       �؇���X�?,            �Q@�      C       D                    4@D�n�3�?             3@        ������������������������       ��<ݚ�?             "@8      ������������������������       ����Q��?             $@      ������������������������       �                     @-      ������������������������       �                     *@,      H       S                 ��Y.@������?J            �\@      I       J                 �?�@(a��䛼?@            @Y@        ������������������������       �                    �E@�       K       R                    �?ܷ��?��?%             M@      L       Q                   �E@ȵHPS!�?!             J@      M       P                   �<@������?            �D@      N       O                 ��) @ףp=
�?             4@      ������������������������       �                     $@�      ������������������������       �z�G�z�?             $@�      ������������������������       �                     5@�       ������������������������       ����|���?             &@      ������������������������       �                     @-      T       U                   @@@և���X�?
             ,@      ������������������������       �؇���X�?             @g      ������������������������       �����X�?             @�       W       X                    �?�FVQ&�?%            �P@        ������������������������       �      �?             @}       Y       Z                 ��T?@ �.�?Ƞ?!             N@       ������������������������       �                    �A@        [       \                   �B@`2U0*��?             9@        ������������������������       �r�q��?             @        ������������������������       �                     3@        �t�bh�h)h,K ��h.��R�(KK]KK��h\�B�        ~@      m@     �d@     �a@     `d@     �D@     �T@      "@      �?      @     �T@      @       @             �R@      @      T@      @@      Q@      ?@      @       @      @      @      @      �?      O@      7@      L@      0@      G@      0@      �?      @     �F@      (@      $@      @      @      @      @             �A@      @      <@      @       @      @      4@              @       @      $@              @      @      (@      �?      @              @      �?      @     �X@      �?      @       @     �W@      �?     �S@      �?      6@      �?      @              2@             �L@      �?      0@      �?      @              "@     �s@      W@     �o@      V@     @P@     �E@      M@       @      $@      @      @       @      @       @      H@      @     �@@              .@      @      @     �A@              @      @      =@      @      8@      @      $@              ,@       @      @     `g@     �F@      U@     �@@     �Q@     �@@     �Q@      :@      @      @      Q@      5@      N@      $@       @      &@       @      @      @      @              @      *@             �Y@      (@     �W@      @     �E@              J@      @      G@      @     �C@       @      2@       @      $@               @       @      5@              @      @      @               @      @      @      �?       @      @      O@      @      @      @     �M@      �?     �A@              8@      �?      @      �?      3@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�
HyhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK	hsK[hth)h,K ��h.��R�(KK[��h{�B�         $                   �'@4�<����?�           @�@                                   �?��̇�?�             s@     �b@                          �1@���|���?3            @S@     �@@������������������������       �      �?              @      9@                           �?8����?.            @Q@     @                          �=@ i���t�?!            �H@     @       
                  s�@؇���X�?            �A@     @       	                 ���@�IєX�?             1@     �X@������������������������       �      �?              @      6@������������������������       �                     "@      0@������������������������       ��<ݚ�?             2@      V@������������������������       �        
             ,@       @                         s�@z�G�z�?             4@      @������������������������       �z�G�z�?             @      8@������������������������       �z�G�z�?	             .@     �F@                          �<@�8(`=��?�            `l@     @                          �;@,I�e���?b            �b@                                 �0@4?,R��?B             [@        ������������������������       �                     *@                                   �?�S����?=            �W@                                  �?z���=��?2            @S@                               ���@��GEI_�?%            �N@        ������������������������       ����Q��?             @        ������������������������       �h�����?!             L@        ������������������������       �     ��?             0@                                  �4@�����H�?             2@        ������������������������       �����X�?             @        ������������������������       �                     &@                                ��) @ �#�Ѵ�?             �E@       ������������������������       �P�Lt�<�?             C@        ������������������������       �z�G�z�?             @                !                 `�X!@���y4F�?1             S@       ������������������������       ��KM�]�?%            �L@3      "       #                    �?�\��N��?             3@       ������������������������       ����!pc�?             &@�       ������������������������       �      �?              @�       %       H                    �?7i����?           �y@       &       /                    �?�q:@Ÿ�?�             m@        '       .                 p"�X@և���X�?             E@       (       )                   �;@`՟�G��?             ?@        ������������������������       ��C��2(�?             &@�       *       +                 ��L@@��Q��?             4@        ������������������������       ������H�?             "@$       ,       -                    E@�eP*L��?             &@        ������������������������       �                     @       ������������������������       �؇���X�?             @-       ������������������������       ��C��2(�?             &@]       0       5                    !@Xf�?s��?u            �g@        1       4                   �C@և���X�?             5@       2       3                    @d}h���?             ,@       ������������������������       �                     $@�       ������������������������       �      �?             @�       ������������������������       �؇���X�?             @�       6       =                 ��D:@��{S�.�?f             e@      7       8                    �?(;L]n�?8            �V@        ������������������������       �"pc�
�?             &@`      9       <                    �?�Fǌ��?0            �S@      :       ;                     @�Ń��̧?             E@      ������������������������       �      �?             @@?      ������������������������       �                     $@I      ������������������������       �                    �B@7      >       E                    �?�2��?.            �S@       ?       D                     @��~R���?$            �O@      @       A                   �G@�\�u��?            �I@      ������������������������       ����"͏�?            �B@�      B       C                   @K@      �?             ,@       ������������������������       �r�q��?             @8       ������������������������       �      �?              @8      ������������������������       ��q�q�?             (@      F       G                 @3#K@      �?
             0@       ������������������������       �                     "@,      ������������������������       �؇���X�?             @�      I       N                     @��!pc�?q             f@       J       K                 ���a@�-.�1a�?J            �^@       ������������������������       �        ?            �Y@v      L       M                 `D�g@ףp=
�?             4@       ������������������������       �      �?              @�      ������������������������       �                     (@�      O       X                    @~|z����?'            �J@      P       Q                    @�e����?            �C@       ������������������������       �                     @�       R       W                 03�7@��.k���?             A@      S       T                    �?����"�?             =@      ������������������������       �X�<ݚ�?             2@%      U       V                   �/@���!pc�?             &@       ������������������������       ����Q��?             @�       ������������������������       �                     @y       ������������������������       �                     @}       Y       Z                    @؇���X�?
             ,@        ������������������������       �r�q��?             @        ������������������������       �      �?              @        �t�bh�h)h,K ��h.��R�(KK[KK��h\�B�        |@     �p@     `n@     �N@     �H@      <@      �?      @      H@      5@      F@      @      >@      @      0@      �?      @      �?      "@              ,@      @      ,@              @      0@      �?      @      @      (@     @h@     �@@     �`@      1@     @W@      .@      *@              T@      .@      P@      *@     �L@      @      @       @      K@       @      @      "@      0@       @      @       @      &@             �D@       @     �B@      �?      @      �?      N@      0@     �I@      @      "@      $@       @      @      �?      @     �i@     `i@     �e@     �L@      8@      2@      ,@      1@      �?      $@      *@      @       @      �?      @      @      @              �?      @      $@      �?     �b@     �C@      "@      (@      @      &@              $@      @      �?      @      �?     �a@      ;@     �U@      @      "@       @     �S@      �?     �D@      �?      ?@      �?      $@             �B@             �K@      8@      D@      7@     �A@      0@      <@      "@      @      @      �?      @      @       @      @      @      .@      �?      "@              @      �?      >@     @b@       @     @^@             �Y@       @      2@       @      @              (@      <@      9@      0@      7@              @      0@      2@      &@      2@       @      $@      @       @      @       @              @      @              (@       @      @      �?      @      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ���]hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKmhth)h,K ��h.��R�(KKm��h{�B@                             �?T�����?�           @�@                                   �?ҳ�wY;�?O            �]@    �S@                           �?��
ц��?6            �S@                               ��>@(���@��?#            �G@                               ���@"pc�
�?            �@@      .@������������������������       �                     @       @       
                   �=@�θ�?             :@              	                 �R,@�����?             3@     0@������������������������       ��q�q�?             (@      @������������������������       �؇���X�?             @      1@������������������������       �                     @      @                         �}S@X�Cc�?
             ,@     �C@������������������������       �r�q��?             @      �?������������������������       �      �?              @       @                            �?��� ��?             ?@                                 �R@R���Q�?             4@      0@������������������������       �      �?              @Z      ������������������������       �                     (@�      ������������������������       ��C��2(�?             &@�                                  @�p ��?            �D@                                 �?      �?             @@       ������������������������       �      �?              @�      ������������������������       �                     8@�      ������������������������       ��<ݚ�?             "@�             V                    �?bN�e�d�?v           ��@                                 !@�繠5�?	           �z@                                  @П[;U��?             =@       ������������������������       �        	             (@                              ��T?@������?	             1@      ������������������������       �                     @(      ������������������������       ����|���?             &@V              '                   �8@�禺f��?�            �x@       !       &                   �4@ ���v��?;            �X@      "       #                     @ףp=
�?              I@       ������������������������       �                      @�       $       %                    �?���H��?             E@       ������������������������       �8�Z$���?             :@v       ������������������������       �      �?             0@j       ������������������������       �                    �H@�       (       5                     �?�w1�|�?�            �r@        )       2                    �?�q�q�?$             K@       *       /                   @>@�(�Tw��?            �C@       +       ,                 ��I/@8�A�0��?             6@        ������������������������       �                     @       -       .                   �J@���Q��?             .@       ������������������������       �      �?              @-       ������������������������       �����X�?             @]       0       1                   �=@�t����?             1@        ������������������������       ��<ݚ�?             "@A       ������������������������       �                      @�       3       4                 03�U@��S���?	             .@       ������������������������       ����Q��?             $@�       ������������������������       ����Q��?             @�       6       U                    �?�}�|���?�            `n@      7       <                   �;@��j���?�            �k@        8       9                     @4�B��?            �B@       ������������������������       �                     $@:      :       ;                   �9@X�<ݚ�?             ;@       ������������������������       �      �?             $@?      ������������������������       �j���� �?	             1@I      =       >                  s�@pb����?u             g@       ������������������������       �                     B@G       ?       T                   �F@�׆���?`            �b@      @       E                   �<@d�;lr�?T            �_@       A       B                 ��@��a�n`�?'             O@       ������������������������       ����Q��?             @�      C       D                    �?l�b�G��?#            �L@        ������������������������       �      �?              @8      ������������������������       ���<D�m�?            �H@      F       M                   @@@      �?-             P@       G       J                 @3�@�q�q�?             ;@       H       I                 �?�@�q�q�?             (@       ������������������������       �z�G�z�?             @�       ������������������������       �և���X�?             @�       K       L                     @������?             .@       ������������������������       �      �?              @�      ������������������������       �����X�?             @�      N       S                    1@��G���?            �B@      O       R                 `fF)@      �?             <@      P       Q                 @3�@�S����?             3@       ������������������������       ��z�G��?             $@�       ������������������������       �                     "@      ������������������������       �X�<ݚ�?             "@-      ������������������������       �                     "@%      ������������������������       �                     7@g      ������������������������       �                     5@�       W       \                     @������?m             e@        X       [                   �:@�"w����?6             S@        Y       Z                   �Y@Pa�	�?            �@@       ������������������������       �                     :@        ������������������������       �؇���X�?             @        ������������������������       �        !            �E@        ]       ^                    .@�û��|�?7             W@        ������������������������       �                     $@        _       b                 ��@�>$�*��?/            �T@        `       a                 ��@@�0�!��?
             1@        ������������������������       �      �?              @        ������������������������       ������H�?             "@        c       j                    �?�4��?%            @P@       d       g                    �?�[�IJ�?            �G@       e       f                   �9@��<b���?             7@        ������������������������       �ףp=
�?             $@        ������������������������       ��	j*D�?             *@        h       i                    �?      �?             8@        ������������������������       �                     @        ������������������������       ��\��N��?             3@        k       l                   �<@�����H�?             2@        ������������������������       �      �?              @        ������������������������       �                     $@        �t�b�`     h�h)h,K ��h.��R�(KKmKK��h\�B�       0|@     Pp@      E@     @S@      B@      E@      @@      .@      ;@      @      @              4@      @      *@      @      @      @      @      �?      @              @      "@      �?      @      @      @      @      ;@      @      1@      @      @              (@      �?      $@      @     �A@      @      <@      @      @              8@       @      @     �y@      g@      v@     @R@      *@      0@              (@      *@      @      @              @      @     0u@     �L@     �W@      @     �F@      @       @             �B@      @      6@      @      .@      �?     �H@             �n@      J@      B@      2@      <@      &@      *@      "@      @              @      "@      �?      @      @       @      .@       @      @       @       @               @      @      @      @       @      @      j@      A@     �g@      A@      9@      (@      $@              .@      (@      @      @      $@      @     `d@      6@      B@             �_@      6@      Z@      6@      L@      @      @       @     �J@      @      @      �?      G@      @      H@      0@      2@      "@      @      @      @      �?      @      @      &@      @      @       @      @       @      >@      @      5@      @      0@      @      @      @      "@              @      @      "@              7@              5@             �L@     �[@      �?     �R@      �?      @@              :@      �?      @             �E@      L@      B@      $@              G@      B@      @      ,@       @      @      �?       @     �E@      6@      ;@      4@      2@      @      "@      �?      "@      @      "@      .@              @      "@      $@      0@       @      @       @      $@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�;hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK
hsKqhth)h,K ��h.��R�(KKq��h{�B@         J                    �?�Qc�!�?�           @�@              ?                 `fFJ@��늓��?)           �|@     @                         ��%@&�~e�?           �y@�y��                            �;@h��� �?�             n@ #y��                              @&<k����?9            @V@     �A@������������������������       �                     @      @                        �Y�@� ��1�?5            �T@      (@       	                    �?      �?             4@     �L@������������������������       ��q�q�?             @      @
                        ��@և���X�?             ,@      J@������������������������       �և���X�?             @        ������������������������       �����X�?             @       @                        ��@��a�n`�?)             O@      @������������������������       �                      @      (@������������������������       ������H�?#             K@      @                          @@@ȨBR��?\             c@     6@                           �?�+�$f��?9            �X@       ������������������������       �z�G�z�?	             .@�                              ��]@�5U��K�?0            �T@                               ���@г�wY;�?             A@       ������������������������       �                     *@n      ������������������������       ����N8�?             5@�                                 ?@؇���X�?            �H@                              ���"@�?�|�?            �B@      ������������������������       �                     @@�      ������������������������       �z�G�z�?             @c      ������������������������       �      �?             (@                                �E@ 7���B�?#             K@      ������������������������       �                     @@�                              pff@�C��2(�?             6@      ������������������������       �        	             ,@V      ������������������������       �      �?              @J      !       $                    @p����?r            �e@       "       #                    @������?             .@      ������������������������       �                     "@�       ������������������������       ��q�q�?             @�       %       6                    �?JN�#:�?e            �c@       &       -                 ��$:@�9�z���?A            @Y@       '       (                   �9@f>�cQ�?$            �N@        ������������������������       �        	             0@�       )       ,                    =@z�G�z�?            �F@        *       +                    �?     ��?             0@        ������������������������       ��q�q�?             @$       ������������������������       �      �?             $@       ������������������������       � 	��p�?             =@       .       5                   �J@��Q��?             D@       /       4                   �>@     ��?             @@       0       1                    �?�t����?             1@        ������������������������       �և���X�?             @A       2       3                 `f�;@ףp=
�?             $@        ������������������������       �                     @�       ������������������������       �z�G�z�?             @�       ������������������������       ���S�ۿ?             .@�       ������������������������       �      �?              @      7       8                    �?@4և���?$             L@        ������������������������       �      �?              @`      9       :                    0@ �q�q�?             H@       ������������������������       �      �?              @;      ;       >                     @�(\����?             D@       <       =                   �A@$�q-�?	             *@       ������������������������       �z�G�z�?             @7      ������������������������       �                      @G       ������������������������       �                     ;@      @       G                   @D@Tt�ó��?"            �H@      A       B                 `f�N@�!���?             A@       ������������������������       �      �?             0@�      C       F                   �;@X�<ݚ�?             2@       D       E                    7@X�<ݚ�?             "@       ������������������������       �      �?             @      ������������������������       ����Q��?             @-      ������������������������       ��q�q�?             "@,      H       I                    �?������?             .@      ������������������������       ��q�q�?             "@�       ������������������������       �r�q��?             @�       K       n                    @�<��S��?�            @o@      L       Y                     @l��N5�?�            �l@      M       V                     �?     �?Q             `@      N       S                    �?      �?-             T@      O       R                    �?���7�?             F@       P       Q                 p��W@�t����?	             1@       ������������������������       �"pc�
�?             &@�       ������������������������       �                     @      ������������������������       �                     ;@-      T       U                 �̴_@�8��8��?             B@      ������������������������       �                     >@g      ������������������������       �      �?             @�       W       X                    6@@��8��?$             H@        ������������������������       ��nkK�?             7@}       ������������������������       �                     9@�       Z       m                   @B@h0�����?=            @Y@       [       \                 ���@j%�*R��?8            @W@        ������������������������       �@4և���?             ,@        ]       f                 ��.@bf@����?1            �S@       ^       _                    �?f�Sc��?             �H@        ������������������������       �                     @        `       a                    �?���Q��?            �F@        ������������������������       ��eP*L��?             &@        b       e                   �9@h+�v:�?             A@       c       d                 pf� @���y4F�?             3@        ������������������������       ��q�q�?             "@        ������������������������       �ףp=
�?             $@        ������������������������       ����Q��?	             .@        g       h                    �?���Q��?             >@        ������������������������       �                     $@        i       l                 ���4@���Q��?             4@       j       k                   �=@և���X�?             ,@        ������������������������       �և���X�?             @        ������������������������       �����X�?             @        ������������������������       �                     @        ������������������������       �                      @        o       p                    �?���N8�?
             5@        ������������������������       �z�G�z�?             $@        ������������������������       ����!pc�?             &@        �t�bh�h)h,K ��h.��R�(KKqKK��h\�B       �{@     �p@      w@     �W@     �u@     �P@     �j@      =@     @R@      0@      @             �P@      0@      $@      $@       @      @       @      @      @      @      @       @      L@      @       @              H@      @     `a@      *@     �U@      &@      (@      @     �R@       @     �@@      �?      *@              4@      �?      E@      @      B@      �?      @@              @      �?      @      @      J@       @      @@              4@       @      ,@              @       @     �`@      C@      @      &@              "@      @       @     @`@      ;@     �S@      7@      J@      "@      0@              B@      "@      "@      @      @       @      @      @      ;@       @      :@      ,@      3@      *@      @      (@      @      @      �?      "@              @      �?      @      ,@      �?      @      �?      J@      @      @       @      G@       @      @      �?     �C@      �?      (@      �?      @      �?       @              ;@              6@      ;@      &@      7@      �?      .@      $@       @      @      @       @       @       @      @      @      @      &@      @      @      @      @      �?     �R@      f@      M@     `e@      @     �^@      @     �R@       @      E@       @      .@       @      "@              @              ;@      @     �@@              >@      @      @      �?     �G@      �?      6@              9@      J@     �H@      F@     �H@      �?      *@     �E@      B@      ?@      2@      @              ;@      2@      @      @      5@      *@      .@      @      @      @      "@      �?      @      "@      (@      2@              $@      (@       @      @       @      @      @       @      @      @               @              0@      @       @       @       @      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ� �thG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKmhth)h,K ��h.��R�(KKm��h{�B@         H                    �?�U��h��?�           @�@              ?                  x#J@@N�Z�=�?           @|@      �                           @�X��)q�?�            0y@      6@                        @3�4@և���X�?             ,@       @������������������������       �                     @      �?������������������������       ��q�q�?             "@      �?       >                 03�>@��C,� �?�            Px@      @       =                   @>@�ڊ��$�?�            `v@      @	       :                   �H@T���D9�?�            �u@      @
       9                 `f�:@4?,R��?�            @t@                                 �:@T�6|���?�            �s@      @                           �?��-�=��?L            @]@     (@                          �9@ܑ-Z���?F            �Z@     @                           �?     ��??             X@       @������������������������       �      �?              @      �?                          �8@`���i��?9             V@     ;@                            @�kb97�?3            @S@       ������������������������       �        	             *@�                              ��Y @      �?*             P@                                �4@�8��8��?             H@                              �?�@�����H�?             ;@      ������������������������       �                     3@�      ������������������������       �      �?              @�                              P��@���N8�?             5@       ������������������������       �z�G�z�?             @�      ������������������������       �        
             0@c      ������������������������       �                     0@      ������������������������       ����!pc�?             &@      ������������������������       �                     &@�      ������������������������       ��z�G��?             $@(             2                   @@@�z����?y            `h@              1                   �?@�9���[�?N            �_@      !       0                   �=@��#:���?F            �[@      "       /                 03�6@Ș����?@             Y@      #       (                    �?��|���?:             V@        $       '                 �R,@�#-���?            �A@       %       &                    �? �Cc}�?             <@        ������������������������       �8�Z$���?
             *@j       ������������������������       ���S�ۿ?
             .@�       ������������������������       �                     @�       )       *                 pb@r�����?!            �J@        ������������������������       �և���X�?             ,@�       +       ,                 ��) @��-�=��?            �C@       ������������������������       �                     5@       -       .                    $@�<ݚ�?             2@        ������������������������       �և���X�?             @-       ������������������������       �                     &@]       ������������������������       ��q�q�?             (@�       ������������������������       �                     $@A       ������������������������       �      �?             0@�       3       8                 ��D:@ ���g=�?+            @Q@       4       5                   �'@`Jj��?'             O@       ������������������������       �                     C@�       6       7                    �?r�q��?             8@      ������������������������       �������?             1@�       ������������������������       �                     @`      ������������������������       �և���X�?             @:      ������������������������       �                     (@;      ;       <                 ���&@ ��WV�?             :@       ������������������������       ��C��2(�?             &@I      ������������������������       �        	             .@7      ������������������������       �      �?              @G       ������������������������       �                     ?@      @       C                    >@և���X�?             �H@       A       B                    �?�eP*L��?             6@       ������������������������       ��z�G��?             $@�      ������������������������       ��q�q�?             (@8       D       E                   �A@�q�q�?             ;@       ������������������������       �                     @      F       G                 03�S@�G�z��?             4@       ������������������������       �����X�?             @,      ������������������������       ���
ц��?             *@�      I       T                     @��&����?�            @p@       J       Q                  "�b@`Ql�R�?X            �a@       K       N                    �? g�yB�?N             `@       L       M                 ��A@��?^�k�?            �A@       ������������������������       �      �?              @�      ������������������������       �                     ;@�      O       P                    �?��K2��?9            �W@      ������������������������       �        !            �M@�      ������������������������       ���?^�k�?            �A@�       R       S                    �?�8��8��?
             (@      ������������������������       �                      @-      ������������������������       �      �?             @%      U       \                    �?@lܯ ��?N            �]@       V       [                    �?�θ�?            �C@       W       X                 Ь* @     ��?             @@       ������������������������       ������?             5@}       Y       Z                    :@���|���?             &@        ������������������������       �z�G�z�?             @        ������������������������       �      �?             @        ������������������������       �և���X�?             @        ]       h                   �>@�z�G��?5             T@       ^       a                   �0@^l��[B�?'             M@        _       `                 �̜6@�C��2(�?	             &@        ������������������������       �      �?             @        ������������������������       �                     @        b       g                 ��Y1@�*/�8V�?            �G@       c       f                    �?^������?            �A@       d       e                   �9@������?             >@       ������������������������       ���s����?             5@        ������������������������       �X�<ݚ�?             "@        ������������������������       �z�G�z�?             @        ������������������������       �                     (@        i       j                   @B@      �?             6@        ������������������������       �ףp=
�?             $@        k       l                 `f(@r�q��?             (@        ������������������������       ����Q��?             @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KKmKK��h\�B�       �z@     �q@     �v@     @V@     `u@     �N@      @       @              @      @      @      u@     �J@     s@     �J@      s@      G@     pq@     �F@     �p@     �F@     @Z@      (@     �X@      "@     �U@      "@      @       @     @T@      @     @R@      @      *@              N@      @      F@      @      8@      @      3@              @      @      4@      �?      @      �?      0@              0@               @      @      &@              @      @     @d@     �@@     @Y@      9@     @W@      1@     �T@      1@     �R@      *@      @@      @      9@      @      &@       @      ,@      �?      @             �E@      $@       @      @     �A@      @      5@              ,@      @      @      @      &@               @      @      $@               @       @     �N@       @      M@      @      C@              4@      @      *@      @      @              @      @      (@              9@      �?      $@      �?      .@              �?      @      ?@              5@      <@      (@      $@      @      @      @      @      "@      2@              @      "@      &@       @      @      @      @      Q@      h@      @     @a@       @     �_@      �?      A@      �?      @              ;@      �?     @W@             �M@      �?      A@      �?      &@               @      �?      @     @P@      K@      "@      >@      @      :@       @      3@      @      @      �?      @      @      @      @      @      L@      8@     �F@      *@      $@      �?      @      �?      @             �A@      (@      7@      (@      6@       @      1@      @      @      @      �?      @      (@              &@      &@      �?      "@      $@       @      @       @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��1hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKshth)h,K ��h.��R�(KKs��h{�B�         0                     @r�����?�           @�@                                  �1@��J�fj�?�            �t@ ��                             �?     ��?             @@        ������������������������       ��<ݚ�?             "@       @                           �?�nkK�?             7@     @������������������������       �                     (@      �?������������������������       ��C��2(�?             &@      @       '                    �?tI��[��?�            �r@     9@	                            �?�0ϔ'6�?l            `f@     @
                        ��$:@Z�K�D��?;            �W@        ������������������������       �                      @                                   �?�&!��?6            �U@     @                          �L@^n����?$             N@     @                        `f�B@H(���o�?            �J@                               ���<@��>4և�?             <@      �?������������������������       ���S���?	             .@      <@                          @C@�θ�?	             *@      ������������������������       �                     @�      ������������������������       �      �?             @�                              `��Z@HP�s��?             9@      ������������������������       �        	             0@n      ������������������������       ��<ݚ�?             "@�      ������������������������       �                     @�                                 �?
j*D>�?             :@       ������������������������       �؇���X�?             @�                              03U@�\��N��?             3@      ������������������������       ��<ݚ�?             "@      ������������������������       ��z�G��?             $@             &                    �?p��@���?1            @U@             !                   �<@�C��2(�?$            �P@                                  �;@r�q��?             >@      ������������������������       �                     2@J      ������������������������       ��q�q�?             (@3      "       %                   �*@������?             B@      #       $                   @D@���7�?             6@       ������������������������       �                     .@�       ������������������������       �؇���X�?             @v       ������������������������       �                     ,@j       ������������������������       �                     3@�       (       -                  "�b@��v$���?P            �^@       )       ,                    �?��wڝ�?G            @[@        *       +                 ��A@h�����?             <@        ������������������������       �      �?              @$       ������������������������       �                     4@       ������������������������       �        6            @T@       .       /                    ;@$�q-�?	             *@        ������������������������       �z�G�z�?             @]       ������������������������       �                      @�       1       ^                    �?���皳�?�            �w@       2       Q                 ��M%@�-x�j�?�            `q@       3       P                 @3�@@mW���?�            �j@       4       O                 �?�@��T��g�?Y            @c@       5       L                   �@������?R            �a@       6       I                 �?$@�v�G���?>            �Y@      7       @                    �?|�M���?3            @U@        8       9                    5@������?            �D@       ������������������������       �����X�?             @:      :       ;                 ���@�IєX�?             A@       ������������������������       �                     *@?      <       ?                   @<@�����?             5@      =       >                    �?      �?             0@       ������������������������       �؇���X�?             @G       ������������������������       �                     "@      ������������������������       �z�G�z�?             @!      A       B                 ��@fP*L��?             F@       ������������������������       �X�<ݚ�?             "@�      C       D                 ���@�#-���?            �A@        ������������������������       �                     (@8      E       F                    7@�LQ�1	�?             7@       ������������������������       �                     $@-      G       H                   �=@�θ�?	             *@      ������������������������       �և���X�?             @�      ������������������������       �                     @�       J       K                   �:@�q�q�?             2@       ������������������������       ������H�?             "@v      ������������������������       �X�<ݚ�?             "@�      M       N                    �?�?�|�?            �B@       ������������������������       �      �?              @�      ������������������������       �                     =@�      ������������������������       �      �?             ,@�      ������������������������       ���S�ۿ?)             N@�       R       S                 ���,@     ��?.             P@       ������������������������       �z�G�z�?             @-      T       [                    �?@�r-��?*            �M@      U       X                    ;@�LQ�1	�?!             G@       V       W                    �?���y4F�?             3@        ������������������������       ��<ݚ�?             "@y       ������������������������       �z�G�z�?             $@}       Y       Z                 03�6@�>����?             ;@       ������������������������       �                     2@        ������������������������       ��<ݚ�?             "@        \       ]                    '@�θ�?	             *@        ������������������������       �և���X�?             @        ������������������������       �                     @        _       l                    �?�7�yHx�?@            @Y@       `       g                 pF @�&�5y�?'             O@        a       d                    �?ܷ��?��?             =@       b       c                 P��@      �?             0@        ������������������������       �z�G�z�?             @        ������������������������       ��C��2(�?             &@        e       f                   �6@$�q-�?             *@        ������������������������       �؇���X�?             @        ������������������������       �                     @        h       k                 pF�-@4���C�?            �@@        i       j                 ��i#@�	j*D�?	             *@       ������������������������       �X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �      �?             4@        m       p                    �?�	j*D�?            �C@        n       o                 ���,@�q�q�?
             .@        ������������������������       �      �?              @        ������������������������       �և���X�?             @        q       r                 �̜6@�8��8��?             8@        ������������������������       �      �?              @        ������������������������       �        
             0@        �t�bh�h)h,K ��h.��R�(KKsKK��h\�B0       �z@      r@      b@     �g@      @      =@       @      @      �?      6@              (@      �?      $@     �a@      d@     `a@      D@      N@      A@       @              J@      A@     �D@      3@      A@      3@      &@      1@       @      @      @      $@              @      @      @      7@       @      0@              @       @      @              &@      .@      �?      @      $@      "@      @       @      @      @     �S@      @      N@      @      9@      @      2@              @      @     �A@      �?      5@      �?      .@              @      �?      ,@              3@               @      ^@      �?      [@      �?      ;@      �?      @              4@             @T@      �?      (@      �?      @               @     �q@     �X@     �m@      E@      g@      =@      `@      9@     �^@      2@     �U@      1@     �R@      &@     �B@      @      @       @      @@       @      *@              3@       @      .@      �?      @      �?      "@              @      �?     �B@      @      @      @      @@      @      (@              4@      @      $@              $@      @      @      @      @              (@      @       @      �?      @      @      B@      �?      @      �?      =@              @      @      L@      @     �I@      *@      �?      @      I@      "@      D@      @      .@      @      @       @       @       @      9@       @      2@              @       @      $@      @      @      @      @              F@     �L@      1@     �F@      @      :@       @      ,@      �?      @      �?      $@      �?      (@      �?      @              @      ,@      3@      "@      @      @      @      @              @      .@      ;@      (@      @      $@      �?      @      @      @      6@       @      @       @      0@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�JIhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK
hsKkhth)h,K ��h.��R�(KKk��h{�B�         Z                 `f~I@������?�           @�@                                   @���[��?m           �@  be use                        ��,)@Nd^����?w            �f@      G@                          �F@�>����?             ;@     (@������������������������       �                     6@       @������������������������       ����Q��?             @      .@                           .@��V��?f            �c@      @������������������������       �                     &@        	                           �?�W�,,T�?^             b@       
                           �?�:���?9            �U@     ^@                            �?�LQ�1	�?,            @Q@     4@                        `f�;@      �?             B@       @                          �H@X�<ݚ�?             "@      9@������������������������       �z�G�z�?             @      @������������������������       �      �?             @       @                        `f�B@PN��T'�?             ;@     �?                        ���=@      �?
             0@       ������������������������       �z�G�z�?             @�      ������������������������       ����!pc�?             &@�      ������������������������       �                     &@w      ������������������������       �                    �@@n                                �?@�X�<ݺ?             2@       ������������������������       �                     $@�      ������������������������       �      �?              @�                                 �?ܷ��?��?%             M@       ������������������������       ����Q��?             @c                                 �?�NW���?!            �J@                                �;@�ʈD��?            �E@       ������������������������       ����Q��?             $@�      ������������������������       �                    �@@(      ������������������������       �                     $@V              ?                    �?�2Ya�Q�?�            �x@      !       $                    $@4?,R��?�             r@       "       #                 ���8@b�2�tk�?
             2@       ������������������������       �                     @�       ������������������������       �                     &@�       %       *                   �5@,sI�v�?�            �p@        &       )                   �0@@�E�x�?            �H@        '       (                    -@$�q-�?             *@        ������������������������       �                      @�       ������������������������       �z�G�z�?             @�       ������������������������       �                     B@�       +       .                    �?8Rq,Y��?�            �k@        ,       -                   �=@��X��?             <@       ������������������������       ��û��|�?             7@       ������������������������       �                     @-       /       8                   @@@(S��C��?u             h@       0       5                   @@��0{9�?V            �a@        1       4                 ��@���?            �D@       2       3                   �:@�r����?             >@        ������������������������       �r�q��?             (@�       ������������������������       ������H�?             2@�       ������������������������       ��eP*L��?             &@�       6       7                 �?�@8EGr��?;             Y@       ������������������������       �                     :@�       ������������������������       ��x
�2�?+            �R@`      9       :                 �?�@ ��WV�?             J@       ������������������������       �                     =@;      ;       >                   �C@���}<S�?             7@      <       =                 �̌!@8�Z$���?	             *@       ������������������������       �����X�?             @7      ������������������������       �                     @G       ������������������������       �                     $@      @       W                   @B@�m��Wv�?D             [@      A       V                     @@��Pl3�?<            @X@      B       Q                    �?�X���?4             V@      C       H                    �?R=6�z�?%            @P@        D       E                   �8@V�a�� �?             =@       ������������������������       ����|���?             &@      F       G                 ���@�����H�?	             2@       ������������������������       �����X�?             @,      ������������������������       �                     &@�      I       J                   �5@*O���?             B@        ������������������������       �      �?              @�       K       N                   �:@      �?             <@      L       M                 P�@�n_Y�K�?
             *@       ������������������������       �                     @�      ������������������������       �����X�?             @�      O       P                 @3�,@�r����?             .@       ������������������������       �؇���X�?             @�      ������������������������       �      �?              @�       R       S                 ��k'@
;&����?             7@       ������������������������       �      �?             @-      T       U                    �?D�n�3�?             3@      ������������������������       ��<ݚ�?             "@g      ������������������������       ����Q��?             $@�       ������������������������       ��<ݚ�?             "@y       X       Y                 0335@�C��2(�?             &@        ������������������������       �z�G�z�?             @�       ������������������������       �                     @        [       h                    �?T��
�?�?P            �`@        \       _                 `�jM@�#}7��?&            �P@        ]       ^                      @�t����?
             1@        ������������������������       �      �?             @        ������������������������       �"pc�
�?             &@        `       c                  D0T@H.�!���?             I@        a       b                    �?P���Q�?             4@        ������������������������       �r�q��?             @        ������������������������       �                     ,@        d       e                 pf�Z@�q�q�?             >@        ������������������������       �      �?              @        f       g                    �?"pc�
�?             6@        ������������������������       ��8��8��?             (@        ������������������������       ��z�G��?             $@        i       j                    �?���7�?*            �P@       ������������������������       �        %             M@        ������������������������       �      �?              @        �t�bh�h)h,K ��h.��R�(KKkKK��h\�B�        |@     `p@     0y@      f@      [@     �R@      9@       @      6@              @       @     �T@     @R@              &@     �T@      O@     @S@      $@      N@      "@      ;@      "@      @      @      �?      @      @      �?      7@      @      (@      @      @      �?       @      @      &@             �@@              1@      �?      $@              @      �?      @      J@       @      @      @     �H@      @     �C@      @      @             �@@              $@     pr@     @Y@      o@      D@      &@      @              @      &@             �m@     �@@      H@      �?      (@      �?       @              @      �?      B@             �g@      @@      3@      "@      ,@      "@      @             @e@      7@      ^@      5@      ?@      $@      :@      @      $@       @      0@       @      @      @     @V@      &@      :@             �O@      &@      I@       @      =@              5@       @      &@       @      @       @      @              $@             �G@     �N@     �B@      N@      >@      M@      3@      G@      @      7@      @      @       @      0@       @      @              &@      *@      7@      @       @      @      5@      @       @              @      @       @       @      *@      �?      @      �?      @      &@      (@      @      �?       @      &@       @      @      @      @      @       @      $@      �?      @      �?      @             �G@     �U@      F@      7@      @      (@      @      @       @      "@     �C@      &@      3@      �?      @      �?      ,@              4@      $@       @      @      2@      @      &@      �?      @      @      @     �O@              M@      @      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��NhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK	hsKOhth)h,K ��h.��R�(KKO��h{�B�                               @Dl���v�?�           @�@                                   �?r�q��?�             u@     �?                           #@�q�q��?t             h@      C@������������������������       �                     $@      @                        ��D:@@S�)�q�?o            �f@                                   4@�zvܰ?0             V@      �?������������������������       ��θ�?             *@     �C@������������������������       �        *            �R@     @Y@	                            �?z�J�??            �W@       
                          �E@�a7���?9            �U@                                 �?@      �?!             I@     "@                          �;@�e����?            �C@      5@                           �?      �?             0@      @������������������������       ��q�q�?             "@      &@������������������������       �և���X�?             @       @������������������������       ���+7��?             7@     �N@������������������������       �"pc�
�?             &@Z                                �L@r�q��?             B@                                 �?�<ݚ�?             ;@       ������������������������       �և���X�?             @w                                �I@R���Q�?             4@      ������������������������       �z�G�z�?	             .@�      ������������������������       �                     @�      ������������������������       �                     "@�      ������������������������       �                      @�                                 @ �q�q�?X             b@       ������������������������       �      �?              @                                 6@ ��ʻ��?T             a@                                 �;@ >�֕�?            �A@       ������������������������       ��<ݚ�?             "@(      ������������������������       �                     :@V      ������������������������       �        @            @Y@J      !       2                    �?�*/�8V�?�            �w@       "       -                    �?nM`����?<             W@      #       &                 P�J@؇>���?(            @P@       $       %                   @<@�MI8d�?            �B@       ������������������������       ��n`���?             ?@v       ������������������������       �                     @j       '       (                    8@X�Cc�?             <@        ������������������������       �      �?              @�       )       ,                   �<@z�G�z�?             4@       *       +                    �?؇���X�?             ,@        ������������������������       �                     @$       ������������������������       �      �?              @       ������������������������       ��q�q�?             @       .       1                 ��.@�q�q�?             ;@       /       0                 Ь* @8�A�0��?             6@       ������������������������       �z�G�z�?
             .@�       ������������������������       �؇���X�?             @A       ������������������������       �                     @�       3       >                    �?����?�            �q@       4       ;                    �?6��m�?�            �i@       5       6                    �?r�q��?y            �f@       ������������������������       �X�If%��?c            �b@      7       8                    1@     ��?             @@        ������������������������       �      �?             @`      9       :                 03S&@@4և���?             <@       ������������������������       ��<ݚ�?             "@;      ������������������������       �                     3@?      <       =                    @`2U0*��?             9@       ������������������������       �r�q��?             @7      ������������������������       �                     3@G       ?       B                   �0@�,�٧��?5            �S@       @       A                    @�r����?             .@       ������������������������       ����Q��?             @�      ������������������������       �                     $@�      C       N                 ���5@     ��?*             P@       D       K                    �?��WV��?!             J@      E       J                    �?      �?             D@      F       G                 ���@�n_Y�K�?             :@       ������������������������       �                     @,      H       I                   �9@�G��l��?             5@      ������������������������       ��	j*D�?             *@�       ������������������������       �      �?              @�       ������������������������       �����X�?             ,@v      L       M                   �*@      �?             (@       ������������������������       �                     @�      ������������������������       �      �?              @�      ������������������������       �        	             (@�      �t�bh�h)h,K ��h.��R�(KKOKK��h\�B�        {@     `q@     @c@     �f@     �b@      F@              $@     �b@      A@     @U@      @      $@      @     �R@             �O@      ?@     �K@      ?@      9@      9@      7@      0@      @      $@      @      @      @      @      1@      @       @      "@      >@      @      5@      @      @      @      1@      @      (@      @      @              "@               @              @     @a@      @      @       @     �`@       @     �@@       @      @              :@             @Y@     �q@      X@      M@      A@     �H@      0@      ?@      @      9@      @      @              2@      $@       @      @      0@      @      (@       @      @              @       @      @       @      "@      2@      "@      *@      @      (@      @      �?              @     �k@      O@     �e@      ?@     �b@      >@     �^@      9@      ;@      @      �?      @      :@       @      @       @      3@              8@      �?      @      �?      3@              H@      ?@      *@       @      @       @      $@             �A@      =@      7@      =@      4@      4@      $@      0@              @      $@      &@      "@      @      �?      @      $@      @      @      "@              @      @      @      (@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ2�3hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKwhth)h,K ��h.��R�(KKw��h{�B�         f                  x#J@l��n�?�           @�@              ?                 `�X.@��*?L�?o           `�@              <                    �?��R[s�?�            �u@      @                           �?���,B�?�            �t@      �?                          �=@n>�X�q�?6             W@     @                        @Q,@� �	��?.            �R@                               ���@$/����?'            @P@     �`@                           �?      �?             <@    @Y@	       
                 ���@�S����?             3@      @������������������������       �                      @      @������������������������       ����!pc�?             &@       @������������������������       �X�<ݚ�?             "@      (@                        ���@V������?            �B@     ?@                        �&B@�q�q�?             >@     @������������������������       ��q�q�?             8@      �?������������������������       ��q�q�?             @       @������������������������       �؇���X�?             @        ������������������������       �                     $@        ������������������������       �                     1@               7                    �?�������?�            �m@                                   @8IMk���?�             i@                                   &@���7�?             F@                                   @�r����?	             .@        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     =@                                  �0@W@e��?d            �c@        ������������������������       �և���X�?             @               6                    �?�r����?`            �b@              /                 @3�@��8���?[            �a@              *                   �>@�㙢�c�?8             W@               )                 �1@pH����?)            �P@       !       &                    :@��G���?            �B@      "       #                   �4@���}<S�?             7@       ������������������������       �                     $@�       $       %                    7@8�Z$���?	             *@       ������������������������       �z�G�z�?             @v       ������������������������       �      �?              @j       '       (                 ���@X�Cc�?             ,@        ������������������������       �r�q��?             @�       ������������������������       �      �?              @�       ������������������������       �                     >@�       +       ,                   @@@��H�}�?             9@        ������������������������       �      �?              @       -       .                   @E@�t����?             1@       ������������������������       �                     &@-       ������������������������       ��q�q�?             @]       0       1                 ��) @�:�]��?#            �I@       ������������������������       �                     <@A       2       5                   �"@�㙢�c�?             7@       3       4                 @Q!@      �?             0@        ������������������������       �      �?             @�       ������������������������       ��8��8��?             (@�       ������������������������       �����X�?             @      ������������������������       �                     @�       8       9                 `fV$@�\��N��?             C@      ������������������������       ��q�q�?             8@:      :       ;                    ?@@4և���?
             ,@       ������������������������       �z�G�z�?             @?      ������������������������       �                     "@I      =       >                    �?D�n�3�?             3@      ������������������������       �X�<ݚ�?             "@G       ������������������������       ����Q��?             $@      @       c                    @����}�?�            �m@      A       X                    �?���m���?�            �j@      B       S                    �?�#DwKd�?P            @^@      C       D                   �9@�������?9            �V@        ������������������������       �                     "@8      E       J                   @<@������?3            @T@       F       G                 ��q1@      �?             @@       ������������������������       �                     @,      H       I                      @X�<ݚ�?             ;@      ������������������������       �D�n�3�?             3@�       ������������������������       �      �?              @�       K       R                   �K@Jm_!'1�?            �H@      L       Q                 ��d;@������?            �B@      M       P                   @D@���y4F�?             3@      N       O                    �?؇���X�?             ,@       ������������������������       �      �?              @�      ������������������������       �r�q��?             @�      ������������������������       ����Q��?             @�       ������������������������       �        	             2@      ������������������������       ��q�q�?             (@-      T       W                     @�4�����?             ?@      U       V                    &@j���� �?             1@       ������������������������       �                     @�       ������������������������       �                     $@y       ������������������������       �d}h���?
             ,@}       Y       \                     @@�҇��?1            �W@       Z       [                    �?`�q�0ܴ?            �G@        ������������������������       �"pc�
�?             &@        ������������������������       �                     B@        ]       b                 ��Y7@��V�I��?            �G@       ^       _                    �?�'�`d�?            �@@        ������������������������       �                     *@        `       a                 03�1@��Q��?             4@        ������������������������       �      �?              @        ������������������������       �      �?             (@        ������������������������       �                     ,@        d       e                    .@���}<S�?             7@       ������������������������       �                     2@        ������������������������       ����Q��?             @        g       r                    �?x�����?M             _@        h       q                    �?ڡR����?!            �H@       i       n                    �?�G��l��?             E@       j       k                   �8@���Q��?             9@        ������������������������       �      �?              @        l       m                    �?��.k���?             1@       ������������������������       ��<ݚ�?             "@        ������������������������       �      �?              @        o       p                     �?j���� �?             1@       ������������������������       ���
ц��?	             *@        ������������������������       �      �?             @        ������������������������       �                     @        s       t                    �?�r����?,            �R@       ������������������������       �        !            �K@        u       v                    @      �?             4@       ������������������������       ����Q��?             .@        ������������������������       �z�G�z�?             @        �t�bh�h)h,K ��h.��R�(KKwKK��h\�Bp       {@     pq@     �x@     @h@     @p@     �V@     �o@     �S@     �M@     �@@      E@     �@@      @@     �@@      5@      @      0@      @       @               @      @      @      @      &@      :@      $@      4@       @      0@       @      @      �?      @      $@              1@              h@      G@     �e@      :@      E@       @      *@       @      @              @       @      =@             �`@      8@      @      @     @`@      4@     �^@      4@      S@      0@      N@      @      >@      @      5@       @      $@              &@       @      @      �?      @      �?      "@      @      @      �?      @      @      >@              0@      "@      �?      @      .@       @      &@              @       @     �G@      @      <@              3@      @      ,@       @      @      �?      &@      �?      @       @      @              2@      4@      1@      @      �?      *@      �?      @              "@       @      &@      @      @      @      @     �`@      Z@     @\@     �Y@     �V@      ?@     @Q@      5@      "@              N@      5@      4@      (@      @              .@      (@      &@       @      @      @      D@      "@     �@@      @      .@      @      (@       @      @      �?      @      �?      @       @      2@              @      @      5@      $@      $@      @              @      $@              &@      @      7@     �Q@       @     �F@       @      "@              B@      5@      :@      @      :@              *@      @      *@      �?      @      @      @      ,@              5@       @      2@              @       @     �C@     @U@      =@      4@      6@      4@      .@      $@      @      �?       @      "@       @      @      @       @      @      $@      @      @      �?      @      @              $@     @P@             �K@      $@      $@      @      "@      @      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJk�ahG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKehth)h,K ��h.��R�(KKe��h{�B@         H                    �?������?�           @�@                                  @�k�+�?7            ~@     �K@                           @���y4F�?             3@     @������������������������       �        	             ,@       @������������������������       �z�G�z�?             @      G@       1                 ��D:@(��?*           �|@                               ��@ą%�E�?�            @v@      @                          �;@ r���?<            �W@      @	       
                 ��@�>����?             ;@       @������������������������       �z�G�z�?             $@      �?������������������������       �                     1@      @������������������������       �        *             Q@      @                         ���!@D�^��?�            Pp@      �?                        �?�@j��>��?O            ``@      4@                          �:@���Ls�?%            @P@      "@                          �5@ 7���B�?             ;@     Z@                          �3@��S�ۿ?	             .@      ������������������������       �                     "@�      ������������������������       �r�q��?             @�      ������������������������       �                     (@w      ������������������������       ��?�'�@�?             C@n                                �E@j�'�=z�?*            �P@                                @@@��$�4��?&            �M@                                �>@      �?             H@                              ��) @��G���?            �B@                                �5@H%u��?             9@       ������������������������       �      �?             @      ������������������������       �                     3@      ������������������������       ��q�q�?	             (@�      ������������������������       ��eP*L��?             &@(      ������������������������       ��C��2(�?             &@V      ������������������������       �և���X�?             @J      !       &                   �4@��a�!��?V            @`@       "       #                     @������?             1@       ������������������������       �r�q��?             @�       $       %                    �?���!pc�?	             &@       ������������������������       �                     @v       ������������������������       ����Q��?             @j       '       *                    �? (��?H            @\@        (       )                 ��$1@��<b���?             7@       ������������������������       ��8��8��?             (@�       ������������������������       ����|���?             &@�       +       ,                   �@@����?�?;            �V@       ������������������������       �        "            �I@       -       0                    �?�7��?            �C@       .       /                   �A@@4և���?             <@        ������������������������       ��q�q�?             @]       ������������������������       �                     6@�       ������������������������       �                     &@A       2       A                    �?�&]�t��?I            �Z@       3       @                     �?      �?1            �R@       4       9                    @@�G��l��?,            �O@        5       8                   �J@      �?             8@       6       7                 0C=@      �?             0@      ������������������������       �z�G�z�?             $@�       ������������������������       �                     @`      ������������������������       �      �?              @:      :       ;                   �;@�n_Y�K�?            �C@       ������������������������       �      �?              @?      <       ?                 ��hU@r֛w���?             ?@      =       >                 `f�B@�LQ�1	�?             7@       ������������������������       ��q�q�?             "@G       ������������������������       �                     ,@      ������������������������       �      �?              @!      ������������������������       ����|���?             &@�      B       G                     �?"pc�
�?            �@@      C       F                 `��`@�����?             3@       D       E                    �?�q�q�?             (@       ������������������������       ��q�q�?             @      ������������������������       �      �?             @-      ������������������������       �؇���X�?             @,      ������������������������       �                     ,@�      I       `                    �?��VT4�?�            �l@       J       O                    �?��9A1�?|            �g@        K       L                     @�����?             E@      ������������������������       �                     =@�      M       N                    .@�	j*D�?	             *@       ������������������������       �                     @�      ������������������������       �և���X�?             @�      P       Y                 `f�$@节>t�?_            �b@       Q       R                    �?      �?             J@        ������������������������       ��t����?             1@      S       T                 ��@���Q��?            �A@       ������������������������       �ףp=
�?             $@%      U       V                   �@z�G�z�?             9@       ������������������������       ����Q��?             @�       W       X                 @3�@R���Q�?             4@        ������������������������       ��<ݚ�?             "@}       ������������������������       ��C��2(�?             &@�       Z       [                     @�^'�ë�?@            @X@       ������������������������       �        ,             Q@        \       _                 03�1@J�8���?             =@       ]       ^                    �?�S����?             3@        ������������������������       �r�q��?             @        ������������������������       �8�Z$���?	             *@        ������������������������       ��z�G��?             $@        a       b                     @��Zy�?            �C@        ������������������������       �@4և���?
             ,@        c       d                 �A7@�J�4�?             9@        ������������������������       �X�<ݚ�?             "@        ������������������������       �        	             0@        �t�bh�h)h,K ��h.��R�(KKeKK��h\�BP        |@     `p@     @x@     �W@      @      .@              ,@      @      �?      x@     �S@      t@      B@     @W@       @      9@       @       @       @      1@              Q@             `l@      A@      [@      7@     �M@      @      :@      �?      ,@      �?      "@              @      �?      (@             �@@      @     �H@      1@      G@      *@      B@      (@      >@      @      6@      @      @      @      3@               @      @      @      @      $@      �?      @      @     �]@      &@      *@      @      @      �?       @      @      @               @      @     �Z@      @      2@      @      &@      �?      @      @      V@       @     �I@             �B@       @      :@       @      @       @      6@              &@              P@     �E@     �B@     �B@     �@@      >@      "@      .@       @      ,@       @       @              @      @      �?      8@      .@      �?      @      7@       @      4@      @      @      @      ,@              @      @      @      @      ;@      @      *@      @      @      @      @       @      @      @      @      �?      ,@              O@      e@      D@     �b@      @      C@              =@      @      "@              @      @      @      B@     @\@      :@      :@      @      (@      5@      ,@      �?      "@      4@      @      @       @      1@      @      @       @      $@      �?      $@     �U@              Q@      $@      3@      @      0@      �?      @       @      &@      @      @      6@      1@      �?      *@      5@      @      @      @      0@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ6ޤhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK
hsKkhth)h,K ��h.��R�(KKk��h{�B�         R                    �? ��ʀ_�?�           @�@              E                 `fFJ@�{���2�?X           X�@     @                            @���<�l�?*           ~@      1@                          @I@ )O7�?]             b@                               `f�B@�Ƀ aA�?M            �]@                                  �?�>���?G             [@     (@                           �?D˩�m��?0            �R@        ������������������������       �      �?             (@      @	                        03�9@t�7��?*             O@     @
                           &@��Y��]�?            �D@      @                           @P���Q�?             4@        ������������������������       �                     @        ������������������������       �$�q-�?             *@      >@������������������������       �                     5@      @                          �E@�G��l��?             5@      @                            �?���Q��?             .@     @������������������������       ��z�G��?             $@Z      ������������������������       ����Q��?             @�      ������������������������       �r�q��?             @�                                @G@г�wY;�?             A@      ������������������������       �                     <@n      ������������������������       �r�q��?             @�      ������������������������       �                     $@�                                  �?���B���?             :@                                @N@������?	             .@       ������������������������       �և���X�?             @c      ������������������������       �      �?              @      ������������������������       ��C��2(�?             &@             0                 ���@Rc����?�            u@              +                    �?��5Е��?R            �`@             *                   �@@(N:!���?A            @Z@              !                    7@R���Q�?0             T@       ������������������������       �`2U0*��?             9@3      "       %                    �?z�G�z�?             �K@       #       $                    �?HP�s��?             9@        ������������������������       �                     @�       ������������������������       ������H�?
             2@v       &       '                 ���@�z�G��?             >@        ������������������������       ��q�q�?             @�       (       )                 pf�@�q�q�?             8@        ������������������������       �                     &@�       ������������������������       ��n_Y�K�?             *@�       ������������������������       �                     9@$       ,       /                 ���@\-��p�?             =@       -       .                 �Y�@��S�ۿ?	             .@        ������������������������       ������H�?             "@-       ������������������������       �                     @]       ������������������������       �d}h���?             ,@�       1       <                    �?< 
2��?{            `i@       2       9                    �?xdQ�m��?`            @d@       3       6                   �3@@��9U��?Q            @a@        4       5                 ��Y @�t����?	             1@        ������������������������       �      �?              @�       ������������������������       �                     "@      7       8                 �?�@���tcH�?H            @^@        ������������������������       �                     C@`      ������������������������       � ,U,?��?1            �T@:      :       ;                   �9@      �?             8@       ������������������������       �      �?              @?      ������������������������       �                     0@I      =       >                    �?#z�i��?            �D@       ������������������������       �      �?             $@G       ?       @                   �7@¦	^_�?             ?@       ������������������������       �                     $@!      A       D                   �>@և���X�?             5@      B       C                 @3�!@X�Cc�?	             ,@      ������������������������       ��q�q�?             "@8       ������������������������       ����Q��?             @8      ������������������������       �և���X�?             @      F       I                    �?����>�?.            �R@       G       H                    �?<���D�?            �@@       ������������������������       �      �?              @�      ������������������������       �                     9@�       J       M                    <@hP�vCu�?            �D@        K       L                   �4@     ��?	             0@       ������������������������       �      �?              @�      ������������������������       �      �?              @�      N       Q                 Ј�U@�q�����?             9@      O       P                    �?�q�q�?	             2@      ������������������������       �                     (@�      ������������������������       �                     @�       ������������������������       �؇���X�?             @      S       \                     @��>���?b            �c@       T       Y                    �?���5��?1            �S@       U       V                    2@�'�=z��?            �@@       ������������������������       �                     .@�       W       X                   �@@�����H�?             2@        ������������������������       �                     "@}       ������������������������       ��<ݚ�?             "@�       Z       [                 ���`@����?�?            �F@       ������������������������       �                    �A@        ������������������������       �ףp=
�?             $@        ]       h                    �?�J�j�?1            �S@       ^       a                 @�+@JJ����?            �G@        _       `                    �?8�Z$���?	             *@        ������������������������       �      �?             @        ������������������������       �                     "@        b       g                    @�!���?             A@       c       d                    $@�5��?             ;@        ������������������������       �                     @        e       f                  �1@z�G�z�?
             4@        ������������������������       �ףp=
�?             $@        ������������������������       ��z�G��?             $@        ������������������������       �                     @        i       j                    @      �?             @@        ������������������������       �؇���X�?             @        ������������������������       �                     9@        �t�b�      h�h)h,K ��h.��R�(KKkKK��h\�B�       �|@     �o@     x@     @e@     �v@      ]@     @V@     �K@      Q@      I@      M@      I@     �L@      1@      @      @     �I@      &@      D@      �?      3@      �?      @              (@      �?      5@              &@      $@      @      "@      @      @      @       @      @      �?      �?     �@@              <@      �?      @      $@              5@      @      &@      @      @      @      @      �?      $@      �?     @q@     �N@     @X@     �B@     @W@      (@      Q@      (@      8@      �?      F@      &@      7@       @      @              0@       @      5@      "@       @      @      3@      @      &@               @      @      9@              @      9@      �?      ,@      �?       @              @      @      &@     `f@      8@      c@      $@     ``@      @      .@       @      @       @      "@              ]@      @      C@             �S@      @      5@      @      @      @      0@              ;@      ,@      @      @      6@      "@      $@              (@      "@      "@      @      @      @      @       @      @      @      4@      K@      @      =@      @      @              9@      0@      9@      @      *@       @      @      �?      @      *@      (@      (@      @      (@                      @      �?      @     @R@      U@      1@     �N@      0@      1@              .@      0@       @      "@              @       @      �?      F@             �A@      �?      "@      L@      7@      9@      6@       @      &@       @       @              "@      7@      &@      0@      &@              @      0@      @      "@      �?      @      @      @              ?@      �?      @      �?      9@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��{hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsK]hth)h,K ��h.��R�(KK]��h{�B@         B                    �?^80�B�?�           @�@              9                  x#J@ӏ�[��?            �|@     @                           @t�Ű�k�?�            �x@      @@                            @      �?             0@      �?������������������������       �                      @     �@@������������������������       �      �?              @      @       .                   �D@ ��P0�?�            �w@     �?       -                    �?�Rez��?�            �s@     (@	                          �0@������?�             r@        
                          �.@�E��ӭ�?	             2@      @������������������������       �      �?              @      9@������������������������       �z�G�z�?             $@      &@                           �?��0k��?�            �p@       @                           @@      �?             @@                                   @`�Q��?             9@                                  �<@���|���?             &@        ������������������������       ��q�q�?             @Z      ������������������������       ����Q��?             @�      ������������������������       �����X�?             ,@�      ������������������������       �                     @w                               ��y @l��\��?�            �m@                              �?�@<���D�?W            �`@                                �;@�8��8��?@             X@       ������������������������       �z�G�z�?             D@�                                  @�h����?!             L@       ������������������������       �                     $@c      ������������������������       ���<b�ƥ?             G@                                �@@�<ݚ�?             B@                              @3�@ �o_��?             9@       ������������������������       ��q�q�?             "@(      ������������������������       �      �?             0@V      ������������������������       ��C��2(�?             &@J      !       "                 `fF)@����?D            �Z@       ������������������������       �                    �B@A      #       ,                     @D��*�4�?/            @Q@       $       +                   �?@,���i�?            �D@       %       *                   �>@      �?             @@       &       '                   �;@�t����?             1@        ������������������������       �                     @�       (       )                   �7@z�G�z�?	             $@       ������������������������       �r�q��?             @�       ������������������������       �      �?             @�       ������������������������       �        	             .@$       ������������������������       ��q�q�?             "@       ������������������������       �                     <@       ������������������������       �        
             8@-       /       0                    �?2L�����?,            @Q@        ������������������������       �r�q��?             @�       1       4                 ��D:@Z���c��?(            �O@       2       3                   @F@ >�֕�?            �A@        ������������������������       �      �?              @�       ������������������������       �                     ;@�       5       8                 �T!@@��>4և�?             <@       6       7                 `f�:@      �?             6@      ������������������������       ���
ц��?             *@�       ������������������������       �X�<ݚ�?             "@`      ������������������������       �                     @:      :       A                    �?$/����?#            @P@      ;       @                     @�E��
��?             J@      <       ?                 �̰f@��6���?             E@      =       >                 Ј�U@�q�q�?            �@@      ������������������������       ��\��N��?             3@G       ������������������������       �؇���X�?             ,@      ������������������������       ������H�?             "@!      ������������������������       �z�G�z�?             $@�      ������������������������       �8�Z$���?             *@�      C       X                 �D�H@ �o_��?�            @o@       D       E                     @�,�:�?_            �d@       ������������������������       �        "             K@      F       W                 ��Y7@�;hѓ��?=            @\@      G       P                   �9@�K��&�?/            �U@      H       I                 ��@X��ʑ��?            �E@       ������������������������       �                      @�       J       M                    �?<=�,S��?            �A@       K       L                   �3@ףp=
�?
             4@       ������������������������       ��q�q�?             @�      ������������������������       �                     ,@�      N       O                    @������?             .@       ������������������������       �؇���X�?             @�      ������������������������       �      �?              @�      Q       V                   �<@��V#�?            �E@       R       U                 ��.@����>�?            �B@      S       T                 �̌@��}*_��?             ;@      ������������������������       �������?             1@%      ������������������������       ����Q��?             $@g      ������������������������       �                     $@�       ������������������������       ��q�q�?             @y       ������������������������       �                     ;@}       Y       \                     �?�}#���?0            �T@       Z       [                    �?�?�|�?+            �R@       ������������������������       �        #             P@        ������������������������       �z�G�z�?             $@        ������������������������       �X�<ݚ�?             "@        �t�bh�h)h,K ��h.��R�(KK]KK��h\�B�       p{@     q@     w@     @W@     u@      N@      @      (@               @      @      @     �t@      H@     `q@      A@     �o@      A@      *@      @      @      @       @       @      n@      =@      8@       @      1@       @      @      @      @       @      @       @      $@      @      @              k@      5@      ]@      0@      V@       @     �@@      @     �K@      �?      $@             �F@      �?      <@       @      2@      @      @      @      (@      @      $@      �?     @Y@      @     �B@              P@      @      B@      @      >@       @      .@       @      @               @       @      @      �?      @      �?      .@              @      @      <@              8@             �K@      ,@      @      �?      I@      *@     �@@       @      @       @      ;@              1@      &@      &@      &@      @      @      @      @      @              @@     �@@      5@      ?@      3@      7@      &@      6@      "@      $@       @      (@       @      �?       @       @      &@       @     �Q@     �f@     �O@      Z@              K@     �O@      I@      B@      I@      6@      5@               @      6@      *@      2@       @      @       @      ,@              @      &@      �?      @      @      @      ,@      =@      $@      ;@      $@      1@      @      *@      @      @              $@      @       @      ;@              @      S@       @      R@              P@       @       @      @      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ?{�hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK
hsK_hth)h,K ��h.��R�(KK_��h{�B�         0                 ��.@�dx<�?�           @�@                                `f#@z����?�            `u@     �?                           �?�����?�            �l@                               �1@(L�\�?�             g@     �@@                        ��@�=C|F�?8            �U@                                 �=@�#-���?-            �Q@     @                           7@�LQ�1	�?             G@       @������������������������       �                     *@      �?	       
                 ��@"pc�
�?            �@@      @������������������������       �և���X�?             @       @������������������������       �ȵHPS!�?             :@      @������������������������       �                     8@      �?������������������������       ��t����?             1@                                  �<@��<D�m�?H            �X@     @������������������������       ����U�?*            �L@      7@                        @3�@������?            �D@      �?                        �?�@z�G�z�?             .@       ������������������������       �ףp=
�?	             $@        ������������������������       ����Q��?             @                                ��i @ ��WV�?             :@                                  @A@�C��2(�?             &@        ������������������������       �r�q��?             @        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       ��q�q�?            �F@               +                   �*@d}h��?F             \@              *                    �?��
ц��?2            �S@              !                   �:@���=�/�?-            @Q@                                  �2@�+$�jP�?             ;@        ������������������������       �      �?              @                                   �'@�}�+r��?             3@       ������������������������       �                     $@        ������������������������       ������H�?             "@3      "       '                    �?և���X�?             E@      #       $                   �@@��s����?             5@        ������������������������       �ףp=
�?             $@�       %       &                 `f�)@���!pc�?	             &@        ������������������������       �z�G�z�?             @j       ������������������������       ��q�q�?             @�       (       )                   `A@���N8�?             5@       ������������������������       �                     ,@�       ������������������������       �؇���X�?             @�       ������������������������       ��<ݚ�?             "@$       ,       -                     @l��\��?             A@        ������������������������       ��q�q�?             @       .       /                   �<@h�����?             <@       ������������������������       �        
             3@]       ������������������������       ������H�?             "@�       1       N                    �?` .�(�?�             w@       2       5                    @ڶ�}��?w            �f@        3       4                   �;@�+e�X�?             9@        ������������������������       ��r����?             .@�       ������������������������       ����Q��?             $@�       6       ?                    �?z\�3�?j            �c@       7       >                     @.�W����?4            �R@       8       =                   �J@@i��M��?,            @P@      9       :                   �>@�n_Y�K�?$             J@       ������������������������       �      �?             8@;      ;       <                 0w�W@�>4և��?             <@      ������������������������       �                     5@I      ������������������������       �����X�?             @7      ������������������������       �$�q-�?             *@G       ������������������������       �      �?             $@      @       K                 ���S@4�{Y���?6            �T@      A       B                    0@$Q�q�?,            �O@       ������������������������       ��q�q�?             @�      C       D                    �?���U�?(            �L@        ������������������������       ������H�?             "@8      E       F                    �?@��8��?!             H@      ������������������������       �                     8@-      G       H                 ��A@ �q�q�?             8@       ������������������������       �                     &@�      I       J                    �?$�q-�?	             *@        ������������������������       �z�G�z�?             @�       ������������������������       �                      @v      L       M                   �B@      �?
             4@       ������������������������       ����|���?             &@�      ������������������������       ��q�q�?             "@�      O       P                    �?�Xbv���?m            `g@       ������������������������       �                     O@�      Q       V                     @@�j���?N            @_@       R       U                   �;@XB���?4            �U@       S       T                   �8@l��\��?             A@      ������������������������       �                     <@%      ������������������������       �      �?             @g      ������������������������       �                    �J@�       W       Z                    �?�d�����?             C@        X       Y                    ;@X�<ݚ�?             2@        ������������������������       ��<ݚ�?             "@�       ������������������������       ��q�q�?             "@        [       ^                    @ףp=
�?             4@       \       ]                   �6@؇���X�?             ,@       ������������������������       �ףp=
�?             $@        ������������������������       �      �?             @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK_KK��h\�B�       �y@     �r@      p@     �U@     �f@     �G@      e@      1@      S@      &@      P@      @      D@      @      *@              ;@      @      @      @      7@      @      8@              (@      @      W@      @     �K@       @     �B@      @      (@      @      "@      �?      @       @      9@      �?      $@      �?      @      �?      @              .@              .@      >@     @R@     �C@      E@      B@      D@      =@      6@      @      @      @      2@      �?      $@               @      �?      2@      8@      1@      @      "@      �?       @      @      @      �?      @       @      �?      4@              ,@      �?      @       @      @      ?@      @      @       @      ;@      �?      3@               @      �?     `c@     �j@      _@     �M@      @      3@       @      *@      @      @     �]@      D@     �H@      :@      F@      5@      @@      4@      "@      .@      7@      @      5@               @      @      (@      �?      @      @     @Q@      ,@     �M@      @      @       @     �K@       @       @      �?     �G@      �?      8@              7@      �?      &@              (@      �?      @      �?       @              $@      $@      @      @      @      @      ?@     �c@              O@      ?@     �W@      @      U@      @      ?@              <@      @      @             �J@      <@      $@      $@       @      @       @      @      @      2@       @      (@       @      "@      �?      @      �?      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��}whG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsK]hth)h,K ��h.��R�(KK]��h{�B@         4                     @�K��?�           @�@               #                  x#J@$/����?�            Pt@     @                           �?�2����?�            �k@     "@                           *@|��"J�?Z            @d@      1@������������������������       �                     @      �?                           �?��t���?V            �c@              
                    �?R�c���?H             `@      =@       	                    =@�\��N��?	             3@       ������������������������       �      �?              @      �?������������������������       ��eP*L��?             &@      4@                          �G@��G�MJ�??            �[@     @                            �?\���(\�?0             T@      �?                          �<@�'�`d�?            �@@     *@������������������������       ��E��ӭ�?             2@      5@                           E@�r����?	             .@        ������������������������       �                     @      ,@������������������������       �      �?              @Z                                 @dP-���?            �G@       ������������������������       �                     "@�                                �<@�KM�]�?             C@       ������������������������       �d}h���?
             ,@n                              `fF)@ �q�q�?             8@       ������������������������       �                     @�      ������������������������       ��IєX�?	             1@�                              `fF:@������?             >@       ������������������������       �@4և���?             ,@c                                �K@     ��?             0@       ������������������������       �؇���X�?             @      ������������������������       ������H�?             "@�      ������������������������       �                     =@(             "                   �;@���#�İ?(            �M@               !                   �7@��S�ۿ?             >@      ������������������������       �                     0@3      ������������������������       �؇���X�?             ,@A      ������������������������       �                     =@�       $       -                    �?>�Q��?B             Z@       %       ,                    �?�GN�z�?(            �P@        &       '                    �?�g�y��?             ?@        ������������������������       ��q�q�?             (@�       (       )                   �?@D�n�3�?             3@        ������������������������       ��q�q�?             @�       *       +                 `fJT@�	j*D�?	             *@       ������������������������       ��<ݚ�?             "@$       ������������������������       �      �?             @       ������������������������       �                    �A@       .       3                 `fmj@�\��N��?             C@       /       0                    �?��X��?             <@        ������������������������       ����Q��?             $@�       1       2                    �?r�q��?             2@       ������������������������       �        
             &@�       ������������������������       �և���X�?             @�       ������������������������       �ףp=
�?             $@�       5       V                 ��Y7@����G��?�            0x@       6       E                    �?f���]�?�            �s@       7       B                 ��.@N֩	%��?4            @V@       8       ?                    �?.}Z*�?)            �Q@      9       >                   @<@z�G�z�?             D@      :       =                    �?������?             >@       ;       <                   �7@b�2�tk�?	             2@       ������������������������       �      �?              @I      ������������������������       ��z�G��?             $@7      ������������������������       ��8��8��?	             (@G       ������������������������       �                     $@      @       A                    9@���@M^�?             ?@       ������������������������       ��q�q�?             (@�      ������������������������       �D�n�3�?
             3@�      C       D                 �=/@r�q��?             2@        ������������������������       �z�G�z�?             $@8      ������������������������       �      �?              @      F       I                 `f#@��m��?�            �l@      G       H                    �?b:�&���?p            �d@      ������������������������       �x�5?,R�?`             b@�      ������������������������       �      �?             6@�       J       O                    �?�4�����?)             O@       K       L                    �?���y4F�?             C@      ������������������������       �                     5@�      M       N                    @@��.k���?             1@      ������������������������       ��q�q�?             (@�      ������������������������       �z�G�z�?             @�      P       S                    0@      �?             8@       Q       R                    �?"pc�
�?             &@        ������������������������       �r�q��?             @      ������������������������       �z�G�z�?             @-      T       U                    �?�θ�?
             *@      ������������������������       �                      @g      ������������������������       ����Q��?             @�       W       X                    �?(N:!���?&            �Q@        ������������������������       ���S���?             .@}       Y       \                    @ �Jj�G�?            �K@       Z       [                    @�g�y��?             ?@        ������������������������       �؇���X�?             @        ������������������������       �                     8@        ������������������������       �                     8@        �t�bh�h)h,K ��h.��R�(KK]KK��h\�B�       @|@     @p@     �d@      d@     �`@     @V@     @`@      @@              @     @`@      <@     @Y@      <@      $@      "@      @      @      @      @     �V@      3@     @Q@      &@      :@      @      *@      @      *@       @      @              @       @     �E@      @      "@              A@      @      &@      @      7@      �?      @              0@      �?      6@       @      *@      �?      "@      @      �?      @       @      �?      =@               @     �L@       @      <@              0@       @      (@              =@     �@@     �Q@      .@     �I@      .@      0@      @       @      &@       @       @      @      "@      @      @       @       @       @             �A@      2@      4@      "@      3@      @      @      @      .@              &@      @      @      "@      �?     �q@      Y@      l@      W@     �G@      E@      F@      ;@      @@       @      6@       @      &@      @      @      @      @      @      &@      �?      $@              (@      3@      @       @       @      &@      @      .@       @       @      �?      @     @f@      I@      a@      >@     @_@      3@      &@      &@      E@      4@      >@       @      5@              "@       @       @      @      �?      @      (@      (@       @      "@      �?      @      �?      @      $@      @       @               @      @      O@       @       @      @      K@      �?      >@      �?      @      �?      8@              8@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�,�hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKshth)h,K ��h.��R�(KKs��h{�B�         P                    �?\H�l�?�           @�@                                   �?
"����?$           �|@      $@                        ���=@��+7��?;             W@       @                        03k:@؇���X�?             <@      *@������������������������       ��z�G��?             $@      @������������������������       ��X�<ݺ?
             2@      �?                           �?     ��?*             P@     @       	                   �>@����S��?&             M@      <@������������������������       �      �?              @     �Q@
                           �?H.�!���?!             I@      @                        �D�J@x�����?            �C@       @                          �=@�X�<ݺ?             2@      @������������������������       �؇���X�?             @      �?������������������������       �                     &@      ;@                           �?�q�q�?             5@     @������������������������       �z�G�z�?             $@      3@������������������������       ��eP*L��?             &@        ������������������������       ����!pc�?             &@        ������������������������       �      �?             @                                   !@�}�J;��?�            �v@                                    @�ՙ/�?             5@        ������������������������       �                     (@                                033>@�����H�?             "@        ������������������������       �                     @        ������������������������       �z�G�z�?             @               M                    �?��0��?�            �u@                                  �?�|��Y��?�            0s@                                `��,@�����?            �H@       ������������������������       ��I�w�"�?             C@        ������������������������       ��C��2(�?             &@               L                    �?�^龆��?�             p@               K                 0��D@\��)��?�            �n@       !       H                    �?X	
bi��?�            @n@      "       #                    �?���\=y�?�             k@       ������������������������       �                     3@�       $       1                     @�C��2(�?            �h@        %       0                   �*@�C��2(�?!            �K@       &       -                   �@@8��8���?             H@       '       (                    @�FVQ&�?            �@@        ������������������������       �                     @�       )       *                    &@@4և���?             <@        ������������������������       �      �?              @�       +       ,                   �;@P���Q�?
             4@       ������������������������       �                     (@       ������������������������       �      �?              @       .       /                   �B@z�G�z�?
             .@        ������������������������       ����Q��?             @]       ������������������������       �ףp=
�?             $@�       ������������������������       �                     @A       2       =                   �;@�C��2(�?^            �a@        3       <                   �8@(��+�?(            �N@       4       7                 ��L@4��?�?!             J@        5       6                  s�@�θ�?	             *@       ������������������������       �r�q��?             @      ������������������������       �����X�?             @�       8       ;                   �3@�7��?            �C@       9       :                 pf� @�r����?             .@      ������������������������       �      �?              @;      ������������������������       �                     @?      ������������������������       �                     8@I      ������������������������       ��q�q�?             "@7      >       C                 �?�@0��P�?6            �T@        ?       B                   �=@ ���J��?            �C@       @       A                 pb@@4և���?
             ,@       ������������������������       �z�G�z�?             @�      ������������������������       �                     "@�      ������������������������       �                     9@8       D       E                 ��y @�ʈD��?            �E@      ������������������������       �H%u��?             9@      F       G                   �<@�X�<ݺ?             2@       ������������������������       �                      @,      ������������������������       �ףp=
�?             $@�      I       J                    +@`2U0*��?             9@        ������������������������       �؇���X�?             @�       ������������������������       �        
             2@v      ������������������������       ����Q��?             @�      ������������������������       �"pc�
�?             &@�      N       O                 �y�/@�?�|�?            �B@       ������������������������       ������H�?             "@�      ������������������������       �                     <@�      Q       d                 ��.@�-��T��?�            �o@        R       [                   �9@���3L�??             [@       S       T                  s�@hP�vCu�?            �D@       ������������������������       �                     "@%      U       Z                   �7@     ��?             @@      V       Y                 �Y5+@��Q��?             4@       W       X                    �?և���X�?             ,@        ������������������������       �      �?             @}       ������������������������       ��z�G��?             $@�       ������������������������       �r�q��?             @        ������������������������       �                     (@        \       c                 �B,@�%o��?(            �P@       ]       `                    �?�������?$             N@        ^       _                 �&B@>���Rp�?             =@       ������������������������       ��t����?	             1@        ������������������������       �r�q��?             (@        a       b                 `f�$@��a�n`�?             ?@        ������������������������       ����|���?             &@        ������������������������       �                     4@        ������������������������       �                     @        e       r                    @��m.	�?[            `b@       f       k                     @������?W            �a@       g       j                   �;@�g�y��?=            @W@        h       i                   �7@ �Cc}�?             <@       ������������������������       �                     2@        ������������������������       ��z�G��?             $@        ������������������������       �        '            @P@        l       m                    �?(���@��?            �G@        ������������������������       �                     .@        n       o                    �?     ��?             @@        ������������������������       �z�G�z�?             .@        p       q                   �8@�t����?             1@       ������������������������       ��<ݚ�?             "@        ������������������������       �      �?              @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KKsKK��h\�B0       �|@     �o@      x@     �Q@      Q@      8@      8@      @      @      @      1@      �?      F@      4@     �D@      1@       @      @     �C@      &@      ?@       @      1@      �?      @      �?      &@              ,@      @       @       @      @      @       @      @      @      @     �s@     �G@       @      *@              (@       @      �?      @              @      �?     `s@      A@      q@     �@@     �C@      $@      =@      "@      $@      �?     `m@      7@     @l@      5@     �k@      3@     �h@      2@      3@             �f@      2@      I@      @     �E@      @      ?@       @      @              :@       @      @      �?      3@      �?      (@              @      �?      (@      @      @       @      "@      �?      @             @`@      *@     �J@       @     �G@      @      $@      @      @      �?      @       @     �B@       @      *@       @      @       @      @              8@              @      @     @S@      @      C@      �?      *@      �?      @      �?      "@              9@             �C@      @      6@      @      1@      �?       @              "@      �?      8@      �?      @      �?      2@              @       @      "@       @      B@      �?       @      �?      <@             �Q@      g@      G@      O@      9@      0@              "@      9@      @      *@      @       @      @      �?      @      @      @      @      �?      (@              5@      G@      ,@      G@      @      6@      @      (@       @      $@      @      8@      @      @              4@      @              9@     �^@      2@     �^@      @     �V@      @      9@              2@      @      @             @P@      .@      @@              .@      .@      1@      @      (@      (@      @      @       @      @      @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�%\hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKghth)h,K ��h.��R�(KKg��h{�B�                             �?^80�B�?�           @�@                                   �?�C��2(�?             &@      "@������������������������       �                     @      D@������������������������       �z�G�z�?             @      3@       H                    �?z�°u�?�           �@    �G@                            �?��!�I�?           |@                                  �9@d��4�o�?;            �W@      $@������������������������       �                     @      5@	                           �?ƈ�VM�?7            @V@      2@
                        �D�G@     ��?             @@        ������������������������       ��<ݚ�?             "@                                   �?\X��t�?             7@     �?                          �?@��.k���?	             1@     @������������������������       �����X�?             @       @������������������������       ��z�G��?             $@        ������������������������       ��q�q�?             @      �?                          �>@�^���U�?$            �L@                                 �<@�����?             3@       ������������������������       �                     @�      ������������������������       �      �?
             (@w                                �B@�I�w�"�?             C@      ������������������������       �      �?             8@�      ������������������������       �        	             ,@�             #                    �?L(ݧa��?�             v@                                   @�θ�?            �C@       ������������������������       �؇���X�?             @c             "                 �&�)@      �?             @@             !                   �=@�q�q�?             8@                              ���@j���� �?             1@       ������������������������       ��q�q�?             @(                                 @@�eP*L��?	             &@      ������������������������       �և���X�?             @J      ������������������������       �      �?             @3      ������������������������       �                     @A      ������������������������       �      �?              @�       $       -                 �?�@�Y���?�            �s@        %       &                 ��@`Ӹ����?8            �V@        ������������������������       �                     C@j       '       (                   �8@$�q-�?             J@        ������������������������       �                     0@�       )       ,                   @@@�����H�?             B@       *       +                   �:@�J�4�?             9@        ������������������������       ��C��2(�?             &@$       ������������������������       �d}h���?             ,@       ������������������������       �                     &@       .       /                    '@���?�             l@        ������������������������       �D�n�3�?             3@]       0       1                 @3�@���z�k�?{            �i@        ������������������������       ��eP*L��?             &@A       2       7                   �9@����H�?t            `h@        3       4                     @ ������?#            �O@        ������������������������       �                     ;@�       5       6                   �2@������?             B@        ������������������������       �                     0@      ������������������������       �P���Q�?             4@�       8       G                   @A@�Ra����?Q            �`@      9       F                    �?�S����?7            �W@      :       E                    �?�=A�F�?.             S@      ;       <                   �;@��$�4��?#            �M@       ������������������������       �      �?              @I      =       B                    ?@��x_F-�?            �I@      >       ?                     @��hJ,�?             A@        ������������������������       ��q�q�?             @      @       A                   �<@ �Cc}�?             <@      ������������������������       ����}<S�?             7@�      ������������������������       �z�G�z�?             @�      C       D                   @@@�t����?	             1@        ������������������������       ����Q��?             @8      ������������������������       �r�q��?             (@      ������������������������       ��t����?             1@-      ������������������������       �        	             3@,      ������������������������       �                    �B@�      I       d                 p�H@����X�?�            �o@       J       K                     @\�$=֢�?w            `h@        ������������������������       �        .            �R@v      L       a                 ��Y7@���?	�?I            @^@      M       P                 ��@�q�q��?<             X@       N       O                    9@��s����?             5@       ������������������������       �                      @�      ������������������������       ��	j*D�?	             *@�      Q       V                  �m#@v�(��O�?-            �R@        R       U                   �;@��a�n`�?             ?@      S       T                   �8@�q�q�?             2@      ������������������������       �"pc�
�?             &@%      ������������������������       �և���X�?             @g      ������������������������       �$�q-�?             *@�       W       Z                   �:@~�4_�g�?             F@        X       Y                 �*@�t����?
             1@        ������������������������       �      �?              @�       ������������������������       ������H�?             "@        [       ^                    �?������?             ;@        \       ]                    �?�n_Y�K�?             *@        ������������������������       �r�q��?             @        ������������������������       �և���X�?             @        _       `                    �?؇���X�?             ,@        ������������������������       �                     $@        ������������������������       �      �?             @        b       c                    @`2U0*��?             9@        ������������������������       �؇���X�?             @        ������������������������       �        	             2@        e       f                    �?0�)AU��?#            �L@       ������������������������       �                    �I@        ������������������������       �r�q��?             @        �t�bh�h)h,K ��h.��R�(KKgKK��h\�Bp       p{@     q@      �?      $@              @      �?      @     `{@     pp@     �v@     �T@      M@     �B@      @              J@     �B@      1@      .@      @       @      $@      *@       @      "@      @       @      @      @       @      @     �A@      6@      @      *@              @      @      @      =@      "@      .@      "@      ,@             @s@      G@      >@      "@      @      �?      8@       @      1@      @      $@      @      @       @      @      @      @      @       @       @      @              @      �?     `q@     �B@     �U@      @      C@              H@      @      0@              @@      @      5@      @      $@      �?      &@      @      &@              h@     �@@       @      &@      g@      6@      @      @     `f@      0@      O@      �?      ;@             �A@      �?      0@              3@      �?     @]@      .@      T@      .@     �N@      .@      G@      *@      @      @     �D@      $@      =@      @      @       @      9@      @      5@       @      @      �?      (@      @       @      @      $@       @      .@       @      3@             �B@              R@     �f@     �Q@      _@             �R@     �Q@      I@     �G@     �H@      @      1@               @      @      "@     �E@      @@      8@      @      (@      @      "@       @      @      @      (@      �?      3@      9@      (@      @      @      @       @      �?      @      4@      @       @      �?      @      @      @       @      (@              $@       @       @      8@      �?      @      �?      2@              �?      L@             �I@      �?      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ2�hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKshth)h,K ��h.��R�(KKs��h{�B�         .                  �#@�Qc�!�?�           @�@               !                    �?6�����?�            �q@Y2	�                              �?���Lͩ�?�             l@     �?                        @� @�C��2(�?�             j@�h��                            @@@�n���k�?r             f@     @                          �?@�?�0�!�?W             a@     G@                        �1@0�v���?S            ``@     @       	                     @L������?.            @R@      @������������������������       �                     $@     �B@
                        ��@�? Da�?(            �O@        ������������������������       ��q�q�?             "@      @                          �:@h�WH��?!             K@      6@������������������������       �        
             5@                                  �=@6YE�t�?            �@@     .@                         s�@�>4և��?             <@      @������������������������       �@4և���?	             ,@      @������������������������       �����X�?
             ,@Z      ������������������������       �                     @�                                �3@XB���?%             M@       ������������������������       �r�q��?             @w                                �<@ pƵHP�?              J@      ������������������������       �                    �C@�      ������������������������       �$�q-�?             *@�      ������������������������       ����Q��?             @�      ������������������������       �                    �D@�                                 ?@     ��?             @@                                �9@��+7��?             7@                                �2@�r����?             .@       ������������������������       �      �?              @�      ������������������������       �                     @(      ������������������������       �      �?              @V      ������������������������       �                     "@J      ������������������������       �      �?             0@3      "       %                    �?�m����?'            �M@       #       $                   �5@�q�q�?             8@        ������������������������       �      �?              @�       ������������������������       �     ��?             0@v       &       '                 ��@���Q��?            �A@        ������������������������       �      �?              @�       (       -                    �?l��
I��?             ;@       )       ,                 `�X!@b�2�tk�?             2@       *       +                   �8@z�G�z�?	             $@       ������������������������       �r�q��?             @$       ������������������������       �      �?             @       ������������������������       �      �?              @       ������������������������       ������H�?             "@-       /       V                     @F��*���?           �z@       0       E                  x#J@���Q��?�            �r@       1       B                    �?�Z����?r            `h@       2       3                   �2@�npº��?\            �b@        ������������������������       �                     &@�       4       ;                    �?և���X�?X            �a@       5       8                    �?�3�E���?@             Z@       6       7                    �?�t����?6            @U@       ������������������������       �և���X�?             @�       ������������������������       �R�}e�.�?1            �S@`      9       :                   �@@�KM�]�?
             3@       ������������������������       ��q�q�?             @;      ������������������������       �                     *@?      <       A                    �?�8��8��?             B@      =       >                    :@ȵHPS!�?             :@       ������������������������       ��<ݚ�?             "@G       ?       @                   �-@�IєX�?             1@      ������������������������       �        	             &@!      ������������������������       �r�q��?             @�      ������������������������       �                     $@�      C       D                    �?��2(&�?             F@        ������������������������       �      �?             (@8      ������������������������       �                     @@      F       I                 p�1N@���{��?B            @Z@       G       H                    �?���7�?             6@       ������������������������       �r�q��?             @�      ������������������������       �                     0@�       J       U                 0U�o@rp��P��?5            �T@       K       P                    �?�M;q��?1            �R@       L       O                   �G@������?             ;@      M       N                    �?�t����?             1@      ������������������������       ��C��2(�?             &@�      ������������������������       �r�q��?             @�      ������������������������       �      �?             $@�      Q       R                  "�b@ �q�q�?             H@       ������������������������       �                     @@      S       T                 `D�c@      �?	             0@       ������������������������       ����Q��?             @%      ������������������������       �                     &@g      ������������������������       �                      @�       W       f                 03c4@     �?^             `@        X       ]                    �?�g�y��?-             O@        Y       Z                    ,@      �?             <@        ������������������������       �                     @        [       \                    �?���}<S�?             7@        ������������������������       ��<ݚ�?             "@        ������������������������       �                     ,@        ^       c                 ��.@�!���?             A@       _       `                    �?      �?             2@        ������������������������       �r�q��?             @        a       b                 ���'@�q�q�?	             (@       ������������������������       �����X�?             @        ������������������������       ����Q��?             @        d       e                    �?      �?             0@        ������������������������       �                     @        ������������������������       �r�q��?             (@        g       j                    �?��2(&�?1            �P@        h       i                    �?�	j*D�?             *@       ������������������������       ��q�q�?             "@        ������������������������       �      �?             @        k       r                 ��p@@0��_��?&            �J@       l       m                    �?��hJ,�?             A@        ������������������������       �                     1@        n       o                    @�t����?             1@        ������������������������       ��q�q�?             @        p       q                 ���7@�C��2(�?	             &@        ������������������������       �r�q��?             @        ������������������������       �                     @        ������������������������       �                     3@        �t�bh�h)h,K ��h.��R�(KKsKK��h\�B0       �{@     �p@      m@     �I@     �i@      5@     �g@      3@     �d@      *@     �^@      *@     @^@      $@     @P@       @      $@             �K@       @      @      @     �H@      @      5@              <@      @      7@      @      *@      �?      $@      @      @              L@       @      @      �?     �I@      �?     �C@              (@      �?       @      @     �D@              :@      @      1@      @      *@       @      @       @      @              @      @      "@              ,@       @      =@      >@       @      0@      @      @      @      *@      5@      ,@       @      @      3@       @      &@      @       @       @      @      �?      @      �?      @      @       @      �?      j@     `k@      ^@     �f@     @X@     �X@     �V@      N@      &@              T@      N@     @S@      ;@      N@      9@      @      @     �L@      5@      1@       @      @       @      *@              @     �@@      @      7@       @      @      �?      0@              &@      �?      @              $@      @      C@      @      @              @@      7@     �T@      �?      5@      �?      @              0@      6@     �N@      6@     �J@      4@      @      .@       @      $@      �?      @      �?      @      @       @      G@              @@       @      ,@       @      @              &@               @     @V@     �C@      @@      >@      5@      @              @      5@       @      @       @      ,@              &@      7@      "@      "@      @      �?      @       @       @      @       @      @       @      ,@              @       @      $@     �L@      "@      "@      @      @      @      @      �?      H@      @      =@      @      1@              (@      @       @      @      $@      �?      @      �?      @              3@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��(.hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsK}hth)h,K ��h.��R�(KK}��h{�B@         4                     @��"{��?�           @�@               !                    �?���Q��?�            `s@     �?                        ���S@�85�r��?            �i@     C@                          @A@��`��?e            �d@     @       
                    �?\X��t�?;             W@     �?                        `fF:@������?#             K@     @������������������������       ��t����?             A@       @       	                   �<@      �?             4@       ������������������������       �     ��?             0@      @������������������������       �      �?             @       @������������������������       �                     C@      �?                        `f�)@ox%�:�?*            @R@     �f@������������������������       ��8��8��?             (@      N@                           G@����5�?#            �N@      5@                           �?� �	��?             9@    �@@                          @D@      �?	             0@     &@������������������������       �                      @Z      ������������������������       �      �?              @�      ������������������������       �                     "@�                                  �?      �?             B@                                �J@���!pc�?             6@       ������������������������       ��n_Y�K�?             *@�      ������������������������       ������H�?             "@�                                �,@d}h���?	             ,@      ������������������������       �                      @�      ������������������������       �      �?             @c                                 �?z�G�z�?             D@                                  �?�����?             3@       ������������������������       �      �?              @�      ������������������������       �                     &@(                                 @B@���N8�?             5@      ������������������������       �                     ,@J      ������������������������       �؇���X�?             @3      "       %                   �8@���N8�?D            @Z@       #       $                 ��D[@h�����?             <@       ������������������������       �                     8@�       ������������������������       �      �?             @v       &       )                 мCG@��cv�?1            @S@        '       (                    �?4���C�?            �@@        ������������������������       �        
             *@�       ������������������������       �P���Q�?             4@�       *       1                  D:T@�GN�z�?             F@       +       0                   �I@ �Cc}�?             <@       ,       /                   @E@R���Q�?             4@       -       .                 ��9L@      �?	             0@       ������������������������       �                     $@-       ������������������������       �r�q��?             @]       ������������������������       �      �?             @�       ������������������������       �                      @A       2       3                    D@     ��?
             0@        ������������������������       �      �?              @�       ������������������������       �      �?              @�       5       b                    �?��5Е��?             y@       6       a                 �T�I@�2����?�            0q@      7       T                    �?�ݰ���?�            �p@       8       9                   �0@�8��8��?�             h@       ������������������������       ��q�q�?             "@:      :       S                   @F@�������?|            �f@      ;       <                 ��@�t����?s            @e@       ������������������������       ����Q��?             @I      =       B                    �?lGts��?o            �d@       >       ?                    ;@r�q��?             B@        ������������������������       �      �?             @      @       A                    �?ףp=
�?             >@      ������������������������       �                     1@�      ������������������������       ��θ�?	             *@�      C       J                 �?�@�ʈD��?V             `@        D       I                 ��L@XB���?(             M@       E       F                   �:@�����H�?             2@       ������������������������       �                     @-      G       H                 pf�@"pc�
�?             &@      ������������������������       �                     @�      ������������������������       ����Q��?             @�       ������������������������       �                     D@�       K       L                 @3�@D��\��?.            �Q@       ������������������������       �X�<ݚ�?             "@�      M       R                 ���#@6uH���?'             O@      N       O                    4@0��_��?             �J@       ������������������������       ����!pc�?             &@�      P       Q                 ���"@���N8�?             E@      ������������������������       �                     @@�       ������������������������       �z�G�z�?             $@      ������������������������       �                     "@-      ������������������������       �        	             *@%      U       \                    5@���@��?,            �R@       V       [                     @p�ݯ��?             C@       W       X                 P�@�q�q�?             8@        ������������������������       �                      @}       Y       Z                 pF�/@      �?             0@        ������������������������       �                     (@        ������������������������       �      �?             @        ������������������������       �        
             ,@        ]       `                  �v6@�X�<ݺ?             B@       ^       _                   �9@�g�y��?             ?@        ������������������������       �؇���X�?             @        ������������������������       �                     8@        ������������������������       �z�G�z�?             @        ������������������������       ��q�q�?             "@        c       z                 ��Y7@�lhM��?M            �_@       d       m                   �7@z�H}��?>            �Z@        e       f                    �?�ʻ����?             A@        ������������������������       ��<ݚ�?             "@        g       l                    �?`�Q��?             9@       h       k                   �5@p�ݯ��?             3@       i       j                 xF4!@��
ц��?
             *@       ������������������������       ��q�q�?             "@        ������������������������       �      �?             @        ������������������������       �r�q��?             @        ������������������������       �r�q��?             @        n       y                   @B@X~�pX��?'            @R@       o       r                   �;@:-�.A�?#            �P@        p       q                   �9@��s����?	             5@        ������������������������       ����Q��?             $@        ������������������������       �                     &@        s       x                    �?�I� �?             G@       t       u                    �?���� �?            �D@       ������������������������       ��LQ�1	�?             7@        v       w                    �?X�<ݚ�?
             2@        ������������������������       �                     @        ������������������������       ��θ�?             *@        ������������������������       �z�G�z�?             @        ������������������������       ��q�q�?             @        {       |                    @P���Q�?             4@       ������������������������       �                     *@        ������������������������       �؇���X�?             @        �t�bh�h)h,K ��h.��R�(KK}KK��h\�B�       �y@     �r@      _@     @g@     �X@     �Z@      W@     @R@      D@      J@      D@      ,@      >@      @      $@      $@      @      "@      @      �?              C@      J@      5@      &@      �?     �D@      4@      ,@      &@      ,@       @       @              @       @              "@      ;@      "@      0@      @       @      @       @      �?      &@      @       @              @      @      @     �@@      @      *@      @       @              &@      �?      4@              ,@      �?      @      9@      T@      �?      ;@              8@      �?      @      8@     �J@      ,@      3@      *@              �?      3@      $@      A@      @      9@      @      1@      �?      .@              $@      �?      @       @       @               @      @      "@      �?      @      @       @     0r@     �[@     �l@     �F@     `l@     �C@      e@      7@      @      @     `d@      4@     �b@      4@      @       @     `b@      2@      >@      @      @      @      ;@      @      1@              $@      @     @]@      (@      L@       @      0@       @      @              "@       @      @              @       @      D@             �N@      $@      @      @     �L@      @      H@      @       @      @      D@       @      @@               @       @      "@              *@              M@      0@      8@      ,@      $@      ,@       @               @      ,@              (@       @       @      ,@              A@       @      >@      �?      @      �?      8@              @      �?      @      @     �N@     �P@      E@     @P@      3@      .@       @      @      1@       @      (@      @      @      @      @      @      �?      @      @      �?      @      �?      7@      I@      3@      H@      @      1@      @      @              &@      .@      ?@      &@      >@      @      4@       @      $@      @              @      $@      @      �?      @       @      3@      �?      *@              @      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJx�+hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKwhth)h,K ��h.��R�(KKw��h{�B�         R                    �?z��Y�)�?�           @�@                                   �?��_	f�?4           �~@                                  @C@(Q����?A            @Y@      @                        03c@F�����?$            �L@     �?                           �?z�J��?            �G@     "@       	                   �>@��6���?             E@      @                          �<@���Q��?             4@     *@������������������������       �����X�?             ,@      ,@������������������������       ��q�q�?             @      8@
                           �?�X����?             6@        ������������������������       ����Q��?             @      1@������������������������       �������?             1@       @������������������������       �                     @       @������������������������       �z�G�z�?             $@      7@                           �?      �?             F@      @                           @@�	j*D�?             :@     @                          �J@և���X�?
             ,@:1	�  ������������������������       ��z�G��?             $@�:1	�  ������������������������       �      �?             @p�$	�  ������������������������       �                     (@�:1	�                             �?r�q��?             2@ :1	�  ������������������������       ����Q��?             @��1	�                            dT@$�q-�?	             *@:1	�  ������������������������       �                      @��1	�  ������������������������       �z�G�z�?             @�:1	�         M                 ��T?@��w"��?�            �x@:1	�                             @0�1a��?�            w@ :1	�  ������������������������       �r�q��?             @�:1	�         D                    @@�𫚛��?�            �v@J��         A                   �*@�F��?�            Pp@:1	�         @                   �>@O�o9%�?�            �j@:1	�          =                    �?�����E�?y            �h@:1	�  !       (                     @���V��?p            �f@       "       #                    @؇���X�?             <@       ������������������������       �                     @�       $       %                   �'@��s����?             5@        ������������������������       �      �?              @v       &       '                   �8@8�Z$���?	             *@       ������������������������       �                      @�       ������������������������       ����Q��?             @�       )       ,                    �?�S����?^             c@        *       +                 ���@      �?             4@        ������������������������       ������H�?             "@$       ������������������������       ����|���?             &@       -       0                 ���@�禺f��?P            �`@        .       /                 P��@��
ц��?             *@        ������������������������       ��q�q�?             @]       ������������������������       �և���X�?             @�       1       :                 ��) @POͳF��?H            �]@       2       3                    �?���F6��?:            �X@        ������������������������       �@4և���?	             ,@�       4       5                   �3@p��@���?1            @U@        ������������������������       �������?             1@�       6       9                   �;@г�wY;�?)             Q@       7       8                   �9@      �?             @@       ������������������������       �                     :@`      ������������������������       ��q�q�?             @:      ������������������������       �                     B@;      ;       <                   �9@�z�G��?             4@      ������������������������       �        
             *@I      ������������������������       �؇���X�?             @7      >       ?                   �5@���y4F�?	             3@       ������������������������       �"pc�
�?             &@      ������������������������       �      �?              @!      ������������������������       �      �?             ,@�      B       C                    +@@��8��?             H@       ������������������������       �؇���X�?             @8       ������������������������       �                    �D@8      E       F                     @г�wY;�?>            �Y@       ������������������������       �                    �G@-      G       H                 �?�@�1�`jg�?%            �K@       ������������������������       �                     @@�      I       L                   `D@�LQ�1	�?             7@       J       K                 pF� @�IєX�?             1@        ������������������������       �r�q��?             @v      ������������������������       �        
             &@�      ������������������������       ��q�q�?             @�      N       Q                    @�q�q�?             8@      O       P                    &@j���� �?             1@       ������������������������       �      �?              @�      ������������������������       ��q�q�?             "@�       ������������������������       �                     @      S       ^                     @�]N���?�            @k@      T       U                    �?`�c�г?N             _@       ������������������������       �                     B@g      V       ]                 03�a@����!p�?8             V@       W       \                   �;@`2U0*��?1            �R@        X       [                    �?ȵHPS!�?             :@        Y       Z                   �7@�θ�?             *@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �        !            �H@        ������������������������       �8�Z$���?             *@        _       f                    �?�ހ��?D            �W@        `       e                    �?�q�q�?             ;@       a       b                   �8@�û��|�?             7@        ������������������������       ��q�q�?             "@        c       d                 ���@d}h���?	             ,@        ������������������������       �      �?             @        ������������������������       �z�G�z�?             $@        ������������������������       �                     @        g       t                    �?�%o��?1            �P@       h       s                    �?\X��t�?"             G@       i       n                 @33"@�Q����?             D@        j       k                 ��@      �?             0@        ������������������������       �      �?             @        l       m                 �?�@�8��8��?             (@        ������������������������       �z�G�z�?             @        ������������������������       �                     @        o       r                    �?      �?             8@        p       q                    4@���!pc�?             &@        ������������������������       �r�q��?             @        ������������������������       ����Q��?             @        ������������������������       ���
ц��?	             *@        ������������������������       �r�q��?             @        u       v                    �?���N8�?             5@        ������������������������       �r�q��?             @        ������������������������       �                     .@        �t�b�@     h�h)h,K ��h.��R�(KKwKK��h\�Bp       �|@     @o@      y@      W@      P@     �B@      ?@      :@      7@      8@      7@      3@       @      (@      @      $@      @       @      .@      @       @      @      *@      @              @       @       @     �@@      &@      2@       @      @       @      @      @      @      �?      (@              .@      @      @       @      (@      �?       @              @      �?      u@     �K@     t@      H@      �?      @      t@     �E@     �k@      D@     �e@     �C@     �d@      @@      c@      <@      8@      @      @              1@      @      @       @      &@       @       @              @       @      `@      8@      .@      @       @      �?      @      @     @\@      3@      @      @      @       @      @      @     �Z@      *@      W@      @      *@      �?     �S@      @      *@      @     �P@       @      >@       @      :@              @       @      B@              ,@      @      *@              �?      @      .@      @      "@       @      @       @      @      @     �G@      �?      @      �?     �D@             �X@      @     �G@              J@      @      @@              4@      @      0@      �?      @      �?      &@              @       @      1@      @      $@      @      @      @      @      @      @              N@     �c@      @     �]@              B@      @     �T@      @      R@      @      7@      @      $@      @      @              @              *@             �H@       @      &@     �K@     �C@      "@      2@      "@      ,@      @      @      @      &@      �?      @       @       @              @      G@      5@      :@      4@      5@      3@      (@      @      �?      @      &@      �?      @      �?      @              "@      .@      @       @      �?      @       @      @      @      @      @      �?      4@      �?      @      �?      .@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJH�SshG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKohth)h,K ��h.��R�(KKo��h{�B�         B                    �?b�`�6��?�           @�@                                   �?�.U֪E�?-           `|@       �                           �?��X��?=             U@                                  �?����X�?9            @S@     �?                          �J@�	j*D�?1            @P@              	                 `f�B@T����1�?+             M@                                ��$:@l��[B��?             =@      @������������������������       �                     @      @@������������������������       ����|���?             6@      @
                        `f&U@д>��C�?             =@      @������������������������       ��}�+r��?             3@      @                          @B@���Q��?             $@      @������������������������       ��q�q�?             @      @������������������������       �      �?             @        ������������������������       �؇���X�?             @        ������������������������       �r�q��?             (@       @������������������������       �����X�?             @              !                 �?�@T}_���?�             w@                                  �;@���۟�?]            `a@                                ��@�r����?            �F@        ������������������������       �X�<ݚ�?             "@                                   �?������?             B@        ������������������������       �r�q��?             @       ������������������������       �                     >@                               ��@`�q�0ܴ?@            �W@                               �Y�@     ��?*             P@                               ���@������?             B@       ������������������������       �                     :@       ������������������������       �ףp=
�?             $@       ������������������������       �                     <@                                  �@ףp=
�?             >@        ������������������������       �      �?              @       ������������������������       �                     6@3      "       7                    �?� ���?�            �l@      #       $                 @3�@H����p�?k            �e@        ������������������������       �      �?              @�       %       6                 0C�E@ĴF���?g            �d@       &       )                    �?@4և���?`            @c@        '       (                    �?      �?             (@        ������������������������       �և���X�?             @�       ������������������������       �                     @�       *       5                   �*@����Q8�?X            �a@       +       ,                 ��) @$�q-�?A             Z@        ������������������������       �                     B@       -       .                    :@�t����?,             Q@        ������������������������       �                     ;@-       /       2                   �=@� ��1�?            �D@        0       1                    $@��S���?             .@       ������������������������       �      �?             $@A       ������������������������       ����Q��?             @�       3       4                 ��Y)@ ��WV�?             :@       ������������������������       �        	             0@�       ������������������������       �ףp=
�?             $@�       ������������������������       �                     C@      ������������������������       ��z�G��?             $@�       8       9                    �?0B��D�?(            �M@       ������������������������       ������H�?             "@:      :       A                     @�:pΈ��?"             I@      ;       <                    *@�q�q�?             8@       ������������������������       �                     @I      =       >                     @�X�<ݺ?             2@       ������������������������       �                      @G       ?       @                   �>@ףp=
�?	             $@       ������������������������       �z�G�z�?             @!      ������������������������       �                     @�      ������������������������       �                     :@�      C       j                    @`�B7��?�             p@       D       M                 `f�$@XeNF���?�            �m@       E       F                    �?��C���?!            �G@       ������������������������       �ҳ�wY;�?             1@-      G       J                   �7@������?             >@       H       I                 �&B@      �?
             (@       ������������������������       �r�q��?             @�       ������������������������       �r�q��?             @�       K       L                   �>@�����H�?
             2@      ������������������������       �                     &@�      ������������������������       �����X�?             @�      N       c                    �?؇���X�?v            �g@      O       ^                   �?@L:�f@�?[            �b@      P       W                     @,�"���?6            @U@      Q       R                     �?`2U0*��?"             I@        ������������������������       �                     4@      S       V                    6@��S�ۿ?             >@      T       U                 `f�)@�r����?             .@       ������������������������       �                     @g      ������������������������       �      �?              @�       ������������������������       �        	             .@y       X       [                    �?">�֕�?            �A@        Y       Z                    �?      �?	             0@        ������������������������       ����Q��?             @        ������������������������       �"pc�
�?             &@        \       ]                    �?p�ݯ��?             3@       ������������������������       ��eP*L��?             &@        ������������������������       �      �?              @        _       `                    G@���7�?%            �P@       ������������������������       �                    �F@        a       b                 ��A@؇���X�?             5@        ������������������������       �      �?              @        ������������������������       �                     *@        d       i                 03�;@p9W��S�?             C@       e       h                    �?�㙢�c�?             7@       f       g                 ��*4@z�G�z�?             .@       ������������������������       ������H�?             "@        ������������������������       ��q�q�?             @        ������������������������       �      �?              @        ������������������������       ���S���?             .@        k       l                  �:@"pc�
�?             6@        ������������������������       �      �?              @        m       n                    @؇���X�?	             ,@       ������������������������       ��q�q�?             @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KKoKK��h\�B�       `|@      p@     �w@     @R@     �L@      ;@     �K@      6@     �F@      4@     �C@      3@      .@      ,@      @               @      ,@      8@      @      2@      �?      @      @      @       @       @       @      @      �?      $@       @       @      @     @t@      G@      `@      $@     �C@      @      @      @     �A@      �?      @      �?      >@             �V@      @     �O@      �?     �A@      �?      :@              "@      �?      <@              ;@      @      @      @      6@             `h@      B@     �b@      5@      �?      @     �b@      ,@     �a@      &@      "@      @      @      @      @             �`@       @      X@       @      B@              N@       @      ;@             �@@       @       @      @      @      @      @       @      9@      �?      0@              "@      �?      C@              @      @      F@      .@      �?       @     �E@      @      1@      @              @      1@      �?       @              "@      �?      @      �?      @              :@             @R@      g@     �K@     �f@      <@      3@      @      &@      6@       @      @      @      �?      @      @      �?      0@       @      &@              @       @      ;@     @d@      0@     �`@      *@      R@       @      H@              4@       @      <@       @      *@              @       @      @              .@      &@      8@      @      (@       @      @       @      "@      @      (@      @      @       @      @      @     �O@             �F@      @      2@      @      @              *@      &@      ;@      @      3@      @      (@      �?       @       @      @      �?      @      @       @      2@      @      @       @      (@       @      @       @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�8�hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKwhth)h,K ��h.��R�(KKw��h{�B�         2                     @�U��h��?�           @�@                                ��\+@��Q�V�?�             t@   

                              @��X��?&             L@      $@������������������������       �                     "@  �                            �?֭��F?�?!            �G@     @       	                    &@��a�n`�?             ?@                                   9@8�Z$���?             *@        ������������������������       ����Q��?             @      @������������������������       �                      @      @
                           C@�X�<ݺ?             2@     @������������������������       �                     $@        ������������������������       �      �?              @      @                        `f�)@      �?             0@        ������������������������       �                     @      .@������������������������       ������H�?             "@      @       +                    �?      �?�            �p@     �?                          �1@�"U����?Z             c@        ������������������������       �                     2@               (                 ��hU@���X�K�?R            �`@                                 �>@���"͏�?E            �[@                                  @=@T����1�?"             M@                                 �A@�3Ea�$�?             G@                                ��";@��Q��?             4@                                  �?��
ц��?	             *@       ������������������������       ��<ݚ�?             "@       ������������������������       �                     @       ������������������������       �                     @                               `fF:@$�q-�?             :@        ������������������������       �                     0@       ������������������������       �z�G�z�?             $@       ������������������������       �r�q��?             (@                #                  x#J@f1r��g�?#            �J@       !       "                   B@�>����?             ;@       ������������������������       ��<ݚ�?             "@A      ������������������������       �                     2@�       $       %                 �D�M@�θ�?             :@        ������������������������       �X�<ݚ�?             "@v       &       '                 �U�R@�IєX�?             1@       ������������������������       �                     (@�       ������������������������       �z�G�z�?             @�       )       *                    �?      �?             8@       ������������������������       �8�Z$���?             *@�       ������������������������       ��C��2(�?             &@$       ,       /                 ���a@�?�|�?J            �[@       -       .                    6@�����?=             W@        ������������������������       �؇���X�?             @-       ������������������������       �        8            @U@]       0       1                    �?�KM�]�?             3@       ������������������������       �                     $@A       ������������������������       ��<ݚ�?             "@�       3       `                    �?      �?�            �x@       4       _                 �T�I@^]X��?�            �q@       5       H                 �?�@H�ՠ&��?�            �p@        6       ?                   �;@�\�)G�?V            �`@       7       >                   �9@     ��?$             H@       8       =                 �1@�p ��?            �D@      9       <                  ��@z�G�z�?             >@      :       ;                    �?      �?             8@       ������������������������       �      �?             @?      ������������������������       �P���Q�?             4@I      ������������������������       �      �?             @7      ������������������������       �        	             &@G       ������������������������       �և���X�?             @      @       G                    �?`��F:u�?2            �U@      A       B                  s�@�:�^���?            �F@       ������������������������       �                     6@�      C       F                    >@�㙢�c�?             7@       D       E                 ��(@������?	             .@      ������������������������       ��<ݚ�?             "@      ������������������������       ��q�q�?             @-      ������������������������       �                      @,      ������������������������       �                     E@�      I       J                 @3�@�h��u�?Y            �`@        ������������������������       �      �?             $@�       K       \                 ��Y7@�0&���?R            @_@      L       M                    ,@�#l��?B            @Y@       ������������������������       �����X�?             @�      N       Y                 03K2@$�3c�s�?<            �W@      O       X                    �?�5U��K�?4            �T@      P       W                   �=@�Z��L��?+            �Q@      Q       V                 ��i @8�Z$���?             J@        R       S                   �3@�+e�X�?             9@       ������������������������       �      �?             @-      T       U                    ;@�S����?
             3@       ������������������������       �                     @g      ������������������������       �      �?             (@�       ������������������������       ��>����?             ;@y       ������������������������       �                     3@}       ������������������������       �        	             (@�       Z       [                 03c4@���!pc�?             &@        ������������������������       �z�G�z�?             @        ������������������������       ��q�q�?             @        ]       ^                    @ �q�q�?             8@        ������������������������       �z�G�z�?             @        ������������������������       �                     3@        ������������������������       ����|���?             &@        a       t                 ���4@.�D�k��?G            �[@       b       q                    �?�0�~�4�?8             V@       c       d                   �0@���e��?)            �P@        ������������������������       �      �?              @        e       p                   �>@�f7�z�?$             M@       f       i                   �7@�n_Y�K�?              J@        g       h                 pff@��.k���?             1@        ������������������������       �z�G�z�?             @        ������������������������       ��q�q�?             (@        j       o                    �?">�֕�?            �A@       k       n                    �?�c�Α�?             =@       l       m                  s�@��<b���?             7@        ������������������������       ��z�G��?             $@        ������������������������       �8�Z$���?             *@        ������������������������       �      �?             @        ������������������������       �      �?             @        ������������������������       ��q�q�?             @        r       s                    .@���!pc�?             6@        ������������������������       �؇���X�?             @        ������������������������       �        
             .@        u       v                    @���}<S�?             7@        ������������������������       ����Q��?             @        ������������������������       �                     2@        �t�bh�h)h,K ��h.��R�(KKwKK��h\�Bp       �z@     �q@      a@     �f@      C@      2@      "@              =@      2@      <@      @      &@       @      @       @       @              1@      �?      $@              @      �?      �?      .@              @      �?       @     �X@     �d@      X@     �L@              2@      X@     �C@      U@      ;@     �C@      3@     �B@      "@      *@      @      @      @       @      @      @              @              8@       @      0@               @       @       @      $@     �F@       @      9@       @      @       @      2@              4@      @      @      @      0@      �?      (@              @      �?      (@      (@       @      &@      $@      �?      @      [@      �?     �V@      �?      @             @U@       @      1@              $@       @      @     `r@     �X@     @n@     �C@     `m@     �A@     �^@      *@     �C@      "@     �A@      @      8@      @      5@      @       @       @      3@      �?      @      @      &@              @      @     �T@      @     �D@      @      6@              3@      @      &@      @      @       @      @       @       @              E@             @\@      6@      @      @      [@      1@     @U@      0@       @      @     �T@      &@     �R@       @     �O@       @      F@       @      3@      @      @      @      0@      @      @              "@      @      9@       @      3@              (@               @      @      @      �?      @       @      7@      �?      @      �?      3@              @      @      J@     �M@      ?@     �L@      9@     �D@      �?      @      8@      A@      4@      @@      "@       @      �?      @       @      @      &@      8@       @      5@      @      2@      @      @       @      &@      @      @      @      @      @       @      @      0@      @      �?              .@      5@       @      @       @      2@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJUehG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKkhth)h,K ��h.��R�(KKk��h{�B�         D                    �?l��n�?�           @�@              /                 ���=@�5*S��?#           0}@     @                           @hau��?�            �v@      @@                        ���3@R���Q�?             4@     �?������������������������       �                     (@        ������������������������       �      �?              @               
                    �?��<���?�            �u@               	                 ��3@&^�)b�?            �E@       ������������������������       �����X�?             <@        ������������������������       �                     .@                                 ��@���79��?�            �r@        ������������������������       �        !             M@                                @3�@h�ʡP��?�            �n@                                �?�@���?2            �T@                                 �4@D|U��@�?)            �P@        ������������������������       �                     &@                                   �?�>4և��?#             L@       ������������������������       �r�q��?             (@�                                �;@"pc�
�?             F@                               �1@�X����?             6@       ������������������������       ��q�q�?             (@n      ������������������������       �                     $@�                                 >@���7�?             6@      ������������������������       �                     .@�      ������������������������       �؇���X�?             @�                                @A@�q�q�?	             .@      ������������������������       �      �?              @      ������������������������       �և���X�?             @             .                 ��D:@ rc����?i            `d@             !                   �3@��Ή�ν?]             b@                                    @     ��?             0@       ������������������������       ������H�?             "@J      ������������������������       �����X�?             @3      "       -                   @A@ �#�Ѵ�?Q             `@      #       &                     @���L��?9            �V@        $       %                   �=@$�q-�?             :@       ������������������������       �                     0@v       ������������������������       �z�G�z�?             $@j       '       (                   �:@����?(            @P@        ������������������������       �                     6@�       )       ,                 `f�'@�ʈD��?            �E@       *       +                   �=@؇���X�?             <@       ������������������������       �@�0�!��?             1@$       ������������������������       ��C��2(�?             &@       ������������������������       �        
             .@       ������������������������       �                     C@-       ������������������������       ��<ݚ�?             2@]       0       C                    @n�ޢ
�?A            @Y@       1       >                   �G@�ҿf���?7            �T@       2       3                 03�>@�U���?*             O@        ������������������������       ��<ݚ�?             "@�       4       7                  x#J@r�z-��?$            �J@        5       6                   �:@�S����?             3@        ������������������������       �      �?             @      ������������������������       �                     *@�       8       =                    >@�ʻ����?             A@      9       <                    �?�q�q�?             8@      :       ;                      @���Q��?	             .@      ������������������������       ����Q��?             @?      ������������������������       ����Q��?             $@I      ������������������������       ������H�?             "@7      ������������������������       �z�G�z�?             $@G       ?       @                   �B@�ՙ/�?             5@       ������������������������       ��<ݚ�?             "@!      A       B                    J@      �?             (@       ������������������������       �����X�?             @�      ������������������������       �z�G�z�?             @8       ������������������������       �        
             2@8      E       j                    @\F~�1�?�            �n@      F       S                     @���GYW�?�            �k@      G       N                   �;@H�Swe�?P            @_@       H       K                   �7@������?            �D@      I       J                    -@h�����?             <@        ������������������������       �؇���X�?             @�       ������������������������       �                     5@v      L       M                   �7@�θ�?
             *@       ������������������������       �      �?             @�      ������������������������       �                     @�      O       R                 ��A@�Ń��̧?3             U@       P       Q                    :@�X�<ݺ?             B@      ������������������������       �                     =@�       ������������������������       �����X�?             @      ������������������������       �                     H@-      T       [                    �?���r
��?D            @X@       U       Z                 ��.@�<ݚ�?            �F@      V       Y                 P��+@����X�?            �A@       W       X                   �5@д>��C�?             =@        ������������������������       ��q�q�?             (@}       ������������������������       ��IєX�?             1@�       ������������������������       �r�q��?             @        ������������������������       �                     $@        \       i                    B@��
ц��?'             J@       ]       h                   �=@�eP*L��?!             F@       ^       e                 `f�%@��+��?            �B@       _       d                   �;@��H�}�?             9@       `       c                 ��,#@�\��N��?             3@       a       b                   �6@�n_Y�K�?             *@       ������������������������       �����X�?             @        ������������������������       �      �?             @        ������������������������       �r�q��?             @        ������������������������       �                     @        f       g                   �:@      �?	             (@       ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �؇���X�?             @        ������������������������       �                      @        ������������������������       ���<b���?             7@        �t�bh�h)h,K ��h.��R�(KKkKK��h\�B�       {@     pq@     0w@      X@     @s@      M@      @      1@              (@      @      @     s@     �D@     �A@       @      4@       @      .@             �p@     �@@      M@             �j@     �@@      O@      4@     �L@      $@      &@              G@      $@      $@       @      B@       @      .@      @      @      @      $@              5@      �?      .@              @      �?      @      $@       @      @      @      @     �b@      *@      a@      "@      *@      @       @      �?      @       @     �^@      @     @U@      @      8@       @      0@               @       @     �N@      @      6@             �C@      @      8@      @      ,@      @      $@      �?      .@              C@              ,@      @     �O@      C@     �F@      C@     �B@      9@       @      @     �A@      2@      0@      @      @      @      *@              3@      .@      1@      @      "@      @      @       @      @      @       @      �?       @       @       @      *@       @      @      @      @       @      @      @      �?      2@              O@     �f@      F@     @f@      @     �]@      @     �B@      �?      ;@      �?      @              5@      @      $@      @      @              @       @     �T@       @      A@              =@       @      @              H@      C@     �M@      $@     �A@      $@      9@      @      8@      @       @      �?      0@      @      �?              $@      <@      8@      4@      8@      3@      2@      0@      "@      $@      "@      @       @       @      @      @      @      @      �?      @              @      "@      @       @              @      �?      @       @              2@      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�)�rhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKOhth)h,K ��h.��R�(KKO��h{�B�         0                    �?��ے@R�?�           @�@                                  �?��Ɛ���?'           p~@                               ��$:@�=��ny�?�            v@                                 @@@X�2{f�?�            0q@     @       
                     @�!�I�*�?{            �g@                                  �(@�S����?             C@        ������������������������       �        	             *@               	                   �;@�+e�X�?             9@       ������������������������       �        
             *@        ������������������������       �      �?             (@        ������������������������       ��h�*$��?a             c@        ������������������������       �        1            @U@                                    @�	j*D�?-            �S@                               �DHC@�G�5��?'            @Q@                                 �<@ҳ�wY;�?             A@                                   �?և���X�?	             ,@        ������������������������       �և���X�?             @Z      ������������������������       �����X�?             @�      ������������������������       �z�G�z�?             4@�                                 �?؇���X�?            �A@                                �@@�C��2(�?             6@      ������������������������       �@4և���?             ,@�      ������������������������       �      �?              @�      ������������������������       ��θ�?             *@�      ������������������������       ��<ݚ�?             "@�                                 @P�~D&�?N            �`@                                 �;@���N8�?             5@      ������������������������       �      �?             0@      ������������������������       �z�G�z�?             @�             +                 ��9L@ ��(��?C            @\@             &                   �9@��O���?2            @U@               %                    �?��G���?            �B@      !       "                     @��Q��?             4@       ������������������������       �z�G�z�?             @A      #       $                    3@���Q��?             .@        ������������������������       ��<ݚ�?             "@�       ������������������������       ��q�q�?             @v       ������������������������       �                     1@j       '       *                     @@��8��?             H@        (       )                   �@@`2U0*��?             9@        ������������������������       �z�G�z�?             @�       ������������������������       �        
             4@�       ������������������������       �                     7@$       ,       /                    �?և���X�?             <@       -       .                    �?�\��N��?             3@        ������������������������       �      �?              @-       ������������������������       ����!pc�?             &@]       ������������������������       ��<ݚ�?             "@�       1       <                     @�1�d��?�             l@       2       3                    &@Xc!J�ƴ?P            �]@        ������������������������       �����X�?             @�       4       7                   �;@�?�|�?L            �[@        5       6                   �8@�}�+r��?             C@       ������������������������       �                    �@@      ������������������������       ����Q��?             @�       8       9                   �H@ �й���?3            @R@      ������������������������       �        '            �K@:      :       ;                 �DD@�X�<ݺ?             2@       ������������������������       �      �?              @?      ������������������������       �                     $@I      =       D                    �?n�tl��?G            �Z@       >       C                 �?�-@0,Tg��?             E@       ?       @                   �0@��>4և�?             <@       ������������������������       �      �?              @!      A       B                 �&B@�G�z��?             4@      ������������������������       ��z�G��?             $@�      ������������������������       ����Q��?             $@8       ������������������������       �                     ,@8      E       L                 �̼6@^��>�b�?.            @P@      F       I                 P��%@�zv�X�?"             F@      G       H                 @3�"@���>4��?             <@      ������������������������       ��ՙ/�?             5@�      ������������������������       �                     @�       J       K                    �?      �?             0@        ������������������������       �      �?              @v      ������������������������       �      �?              @�      M       N                    #@���N8�?             5@       ������������������������       �؇���X�?             @�      ������������������������       �                     ,@�      �t�bh�h)h,K ��h.��R�(KKOKK��h\�B�       �|@     �o@     `y@     @T@     @s@     �F@     �o@      5@      e@      5@      @@      @      *@              3@      @      *@              @      @      a@      .@     @U@              K@      8@      J@      1@      6@      (@      @       @      @      @       @      @      0@      @      >@      @      4@       @      *@      �?      @      �?      $@      @       @      @     �X@      B@      @      0@      �?      .@      @      �?     @W@      4@     @S@       @      >@      @      *@      @      @      �?      "@      @      @       @       @      @      1@             �G@      �?      8@      �?      @      �?      4@              7@              0@      (@      "@      $@      �?      @       @      @      @       @     �J@     �e@      @     @\@       @      @      @      [@       @      B@             �@@       @      @      �?      R@             �K@      �?      1@      �?      @              $@      H@     �M@      &@      ?@      &@      1@       @      @      "@      &@      @      @      @      @              ,@     �B@      <@      1@      ;@      .@      *@       @      *@      @               @      ,@      �?      @      �?      @      4@      �?      @      �?      ,@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJX"4qhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK
hsKahth)h,K ��h.��R�(KKa��h{�B@         &                 ��%@�3�n��?�           @�@               	                    �?܈=�Z��?�            �q@      @                           �?�q�q�?/            @Q@     &@������������������������       ���p\�?            �D@                                ���@����X�?             <@                                   �?z�G�z�?	             .@        ������������������������       �                      @        ������������������������       �և���X�?             @       ������������������������       ��n_Y�K�?	             *@        
                          �4@0��xX��?�            @k@                                  �3@������?            �D@                               �?�@      �?             @@       ������������������������       �                     4@       ������������������������       �r�q��?             (@       ������������������������       �                     "@               #                    �?@�r-��?w             f@                                 �;@�	L �F�?e            `c@                                ���@     ��?             @@        ������������������������       ��q�q�?             @        ������������������������       �ȵHPS!�?             :@                                �?�@4Qi0���?N            �^@                               ��@�g�y��?)             O@        ������������������������       �                     <@                                  �@�IєX�?             A@        ������������������������       �"pc�
�?             &@        ������������������������       �                     7@                                @3�@f>�cQ�?%            �N@        ������������������������       �����X�?             @               "                   @@@�>����?             K@              !                 ���"@�t����?             A@                                  �=@P���Q�?             4@       ������������������������       �        	             *@        ������������������������       �؇���X�?             @3      ������������������������       �d}h���?             ,@A      ������������������������       �                     4@�       $       %                 P�@8�A�0��?             6@        ������������������������       ��q�q�?             @v       ������������������������       �     ��?             0@j       '       N                    �?*�V����?           �z@       (       =                     �?�P�����?�            �o@        )       2                   �>@��k��?<            �Z@        *       1                 ���=@�ՙ/�?             E@       +       0                   @K@��S���?             >@       ,       /                 ��";@���!pc�?             6@       -       .                 03k:@      �?             0@        ������������������������       �����X�?             @-       ������������������������       �                     "@]       ������������������������       ��q�q�?             @�       ������������������������       �                      @A       ������������������������       �r�q��?             (@�       3       8                 Ј�U@     ��?%             P@       4       5                   �;@R���Q�?             D@        ������������������������       ����Q��?             @�       6       7                 �K@b�h�d.�?            �A@      ������������������������       �������?
             1@�       ������������������������       ������H�?	             2@`      9       <                    �?r�q��?             8@      :       ;                   �D@�θ�?             *@       ������������������������       �؇���X�?             @?      ������������������������       ��q�q�?             @I      ������������������������       ����!pc�?             &@7      >       A                    @��[.K�?\            @b@        ?       @                    @�z�G��?             4@      ������������������������       �                     (@!      ������������������������       �      �?              @�      B       K                    �?|�(��?P            �_@      C       J                 0��D@0)RH'�?+            @Q@       D       I                 ��q1@ףp=
�?&             N@      E       H                 ���+@HP�s��?             I@      F       G                   �;@�����?             E@       ������������������������       �                     *@,      ������������������������       �\-��p�?             =@�      ������������������������       �                      @�       ������������������������       �z�G�z�?             $@�       ������������������������       �X�<ݚ�?             "@v      L       M                 ��Y/@���U�?%            �L@       ������������������������       ��q�q�?             @�      ������������������������       �        !            �I@�      O       `                    @���PL6�?k            �e@      P       [                 039@1�	�?e            �d@       Q       Z                   �E@����O��?(            �Q@       R       Y                    7@�w��@�?$            �O@      S       V                    �?���c���?              J@      T       U                    �?Pa�	�?            �@@      ������������������������       �                     6@g      ������������������������       ��C��2(�?             &@�       W       X                  �2@�����?             3@       ������������������������       ��eP*L��?             &@}       ������������������������       �      �?              @�       ������������������������       �"pc�
�?             &@        ������������������������       �      �?              @        \       _                     @heu+��?=            �W@       ]       ^                 03�a@�x�E~�?8            @V@       ������������������������       �        /             R@        ������������������������       ��t����?	             1@        ������������������������       �                     @        ������������������������       �      �?              @        �t�bh�h)h,K ��h.��R�(KKaKK��h\�B       �{@     �p@     `m@      J@      G@      7@      C@      @       @      4@      @      (@               @      @      @      @       @     �g@      =@     �C@       @      >@       @      4@              $@       @      "@             �b@      ;@      a@      2@      9@      @       @      @      7@      @      \@      &@      N@       @      <@              @@       @      "@       @      7@              J@      "@       @      @      I@      @      >@      @      3@      �?      *@              @      �?      &@      @      4@              *@      "@       @      @      &@      @     `j@     �j@      f@     �R@      M@      H@      0@      :@      ,@      0@      @      0@       @      ,@       @      @              "@      @       @       @               @      $@      E@      6@      ?@      "@       @      @      =@      @      *@      @      0@       @      &@      *@      @      $@      �?      @       @      @       @      @     �]@      ;@      @      ,@              (@      @       @     @\@      *@      M@      &@      K@      @      G@      @      C@      @      *@              9@      @       @               @       @      @      @     �K@       @      @       @     �I@              A@     `a@      <@      a@      5@      I@      0@     �G@      @     �F@      �?      @@              6@      �?      $@      @      *@      @      @      �?      @      "@       @      @      @      @     �U@       @     �U@              R@       @      .@      @              @       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ;�3whG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKyhth)h,K ��h.��R�(KKy��h{�B@         T                    �?(����7�?�           @�@                                  �?|(:�ޞ�?           p|@      1@                          @@.Lj���?.             Q@      �?������������������������       �      �?	             0@       @                           �?
j*D>�?%             J@     @                           �?���Q��?             D@     @                         �}S@�q�q�?             ;@     .@                          �<@���Q��?             4@     @	       
                     �?�	j*D�?
             *@       @������������������������       �և���X�?             @      �?������������������������       �r�q��?             @      (@������������������������       �և���X�?             @       @������������������������       �؇���X�?             @      [@                        �D�C@��
ц��?	             *@      R@������������������������       �և���X�?             @      $@������������������������       ��q�q�?             @      @                           6@      �?             (@       ������������������������       �                     @�      ������������������������       �      �?              @�                                 @�T|n�q�?�            0x@                                   @�㙢�c�?
             7@       ������������������������       �                     &@�      ������������������������       ��q�q�?             (@�             %                     �?Ĝ�oV4�?�            �v@                                �T!@@j�g�y�?&             O@                               `fF<@��
ц��?             :@                              ��$:@�E��ӭ�?             2@       ������������������������       �                     @                                �J@�q�q�?             (@       ������������������������       �����X�?             @(      ������������������������       �                     @V      ������������������������       �      �?              @J      !       "                   �;@�8��8��?             B@       ������������������������       �"pc�
�?             &@A      #       $                    �?`2U0*��?             9@       ������������������������       �                     3@�       ������������������������       �r�q��?             @v       &       M                    �?(+ �8�?�            �r@       '       L                 0�_F@��O���?�            �l@       (       )                   �2@�����?�            �k@        ������������������������       �                     7@�       *       G                 `f�&@̧�*�?�            �h@       +       D                   �E@�r����?g            �b@       ,       C                   �C@���H��?]            �`@       -       B                 ���!@(��+�?X            �^@       .       A                 ��) @����X��?M            @Z@       /       <                 �?�@ ���3�?I            �X@       0       ;                 �1@�qM�R��?5            �P@       1       :                    =@��E�B��?"            �G@       2       5                    7@@�0�!��?             A@        3       4                   �5@$�q-�?	             *@       ������������������������       �؇���X�?             @�       ������������������������       �                     @�       6       7                   �;@���N8�?             5@       ������������������������       ����Q��?             @�       8       9                 03�@     ��?             0@       ������������������������       �                     @:      ������������������������       ����!pc�?             &@;      ������������������������       �                     *@?      ������������������������       �                     4@I      =       >                 @3�@     ��?             @@       ������������������������       �X�Cc�?             ,@G       ?       @                    ;@�����H�?             2@       ������������������������       ����Q��?             @!      ������������������������       �        	             *@�      ������������������������       �      �?             @�      ������������������������       �                     1@8       ������������������������       �                     &@8      E       F                 pff@������?
             1@       ������������������������       �                     $@-      ������������������������       �և���X�?             @,      H       K                   �*@@�E�x�?            �H@       I       J                   �@@�nkK�?             7@       ������������������������       �        	             ,@�       ������������������������       ������H�?             "@v      ������������������������       �                     :@�      ������������������������       �؇���X�?             @�      N       O                    !@��pBI�?)            @R@       ������������������������       �z�G�z�?             @�      P       Q                    ?@ ��ʻ��?%             Q@      ������������������������       �                     J@�       R       S                   �A@      �?             0@       ������������������������       �      �?             @-      ������������������������       �                     (@%      U       ^                   �5@�\T����?�            p@       V       ]                 ���I@X�<ݚ�?'            �O@       W       X                     @D7�J��?!            �K@        ������������������������       �        	             &@}       Y       Z                 �*@���|���?             F@       ������������������������       �\X��t�?             7@        [       \                    �?؇���X�?             5@        ������������������������       ��z�G��?             $@        ������������������������       �                     &@        ������������������������       �                      @        _       r                    �?���*�?            @h@       `       k                    �?Z�J�p�?k            �d@       a       b                    �?���c���?E             Z@        ������������������������       �г�wY;�?             A@        c       f                   �9@z��R[�?,            �Q@        d       e                     @���|���?	             &@        ������������������������       �z�G�z�?             @        ������������������������       �      �?             @        g       h                     @@�r-��?#            �M@       ������������������������       �                    �C@        i       j                 `�X!@�G�z��?             4@       ������������������������       ��q�q�?             (@        ������������������������       �      �?              @        l       o                     @�&�5y�?&             O@       m       n                    :@P���Q�?             D@        ������������������������       ��<ݚ�?             "@        ������������������������       �                     ?@        p       q                    �?�X����?             6@        ������������������������       ��q�q�?             (@        ������������������������       �z�G�z�?             $@        s       t                   �8@և���X�?             <@        ������������������������       �                     $@        u       v                     @�q�q�?             2@        ������������������������       ����Q��?             @        w       x                    �?�θ�?
             *@        ������������������������       �և���X�?             @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KKyKK��h\�B�       �{@      q@     w@     �U@     �F@      7@      .@      �?      >@      6@      8@      0@      2@      "@      (@       @      "@      @      @      @      @      �?      @      @      @      �?      @      @      @      @       @      @      @      @              @      @       @     @t@     �O@      @      3@              &@      @       @      t@      F@     �G@      .@      ,@      (@      *@      @      @              @      @       @      @      @              �?      @     �@@      @      "@       @      8@      �?      3@              @      �?     q@      =@     @i@      ;@      i@      5@      7@             @f@      5@     @`@      4@     @]@      0@     �Z@      0@     @V@      0@     �U@      *@     �N@      @     �D@      @      <@      @      (@      �?      @      �?      @              0@      @      @       @      *@      @      @               @      @      *@              4@              9@      @      "@      @      0@       @      @       @      *@              @      @      1@              &@              *@      @      $@              @      @      H@      �?      6@      �?      ,@               @      �?      :@              �?      @     �Q@       @      @      �?     �P@      �?      J@              .@      �?      @      �?      (@             �Q@     @g@      <@     �A@      <@      ;@              &@      <@      0@      $@      *@      2@      @      @      @      &@                       @     �E@     �b@      ?@     �`@      ,@     �V@      �?     �@@      *@     �L@      @      @      �?      @      @      @      "@      I@             �C@      "@      &@      @      @       @      @      1@     �F@       @      C@       @      @              ?@      .@      @      @      @       @       @      (@      0@              $@      (@      @       @      @      $@      @      @      @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�3hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKihth)h,K ��h.��R�(KKi��h{�B@         H                    �?(����7�?�           @�@                                  @F.< ?�?&           �|@                                   @���N8�?             5@     *@������������������������       �        
             .@      @������������������������       �r�q��?             @     @                           �?��m.	�?           �{@      @                           5@��Q:��?)            �M@      .@������������������������       �����X�?             @     @	       
                 ���<@θ	j*�?$             J@      @������������������������       ��+e�X�?             9@      �?                           �?�5��?             ;@     (@                          �A@���|���?             6@       @������������������������       ����Q��?             @      [@                         "�e@�t����?             1@      R@������������������������       �"pc�
�?             &@      $@������������������������       �      �?             @      @������������������������       ����Q��?             @Z             9                 ��D:@x�v�#��?�            �w@             &                 @3�@��P��i�?�            �q@              %                   �E@F�4�Dj�?M            �]@             "                    �?�L"��?I            �Z@                                  @Df/��?A            �W@       ������������������������       �                     $@�                                �4@0,Tg��?9             U@       ������������������������       �        	             ,@�             !                 �?�@z��R[�?0            �Q@                                �;@Xny��?,            �N@                               ��L@     ��?             0@      ������������������������       ��eP*L��?             &@�      ������������������������       �                     @(                                  �?`Ӹ����?             �F@       ������������������������       �z�G�z�?             $@J      ������������������������       �                    �A@3      ������������������������       ��q�q�?             "@A      #       $                   �7@�	j*D�?             *@        ������������������������       �      �?              @�       ������������������������       �z�G�z�?             @v       ������������������������       ��eP*L��?             &@j       '       2                     @�@�?g            `d@        (       1                    �?t�e�í�?+            �P@       )       0                    F@�.ߴ#�?'            �N@       *       -                   �@@      �?             H@       +       ,                    &@Pa�	�?            �@@        ������������������������       �ףp=
�?             $@       ������������������������       �                     7@       .       /                   �A@�r����?	             .@        ������������������������       �r�q��?             @]       ������������������������       ������H�?             "@�       ������������������������       �                     *@A       ������������������������       ��q�q�?             @�       3       8                    �?      �?<             X@       4       7                 `f�'@p�C��?8            �V@       5       6                 ���"@�&=�w��?"            �J@       ������������������������       �@��8��?             H@      ������������������������       �z�G�z�?             @�       ������������������������       �                     C@`      ������������������������       �z�G�z�?             @:      :       E                    �?�9�z���?;            @Y@      ;       D                     @��Q��?%             N@      <       ?                   �>@�t����?            �I@       =       >                   @=@�G��l��?             5@      ������������������������       ����Q��?	             .@G       ������������������������       �r�q��?             @      @       C                    D@�r����?             >@      A       B                   @K@"pc�
�?             6@       ������������������������       ��C��2(�?             &@�      ������������������������       ����!pc�?             &@8       ������������������������       �                      @8      ������������������������       ��q�q�?             "@      F       G                    !@������?            �D@       ������������������������       �r�q��?             (@,      ������������������������       �                     =@�      I       V                   �5@[z4Փ�?�            @o@        J       K                     @�):u��?+            @S@        ������������������������       �                     7@v      L       M                    �?�q�q�?             K@       ������������������������       �                     @�      N       S                    �?      �?             H@      O       P                  s�@�n_Y�K�?             :@       ������������������������       �      �?             (@�      Q       R                 @� @@4և���?	             ,@        ������������������������       �z�G�z�?             @      ������������������������       �                     "@-      T       U                    @�C��2(�?
             6@       ������������������������       ��<ݚ�?             "@g      ������������������������       �                     *@�       W       X                 `f�$@�%�@>��?j            �e@        ������������������������       �hP�vCu�?            �D@}       Y       d                     @��U�=��?R            �`@       Z       _                   �;@�]��??            �Y@        [       ^                 83�`@     ��?             @@       \       ]                    �? ��WV�?             :@       ������������������������       ��C��2(�?             &@        ������������������������       �                     .@        ������������������������       ��q�q�?             @        `       a                   �H@ ��PUp�?.            �Q@       ������������������������       �        $            �K@        b       c                    �?      �?
             0@        ������������������������       �r�q��?             @        ������������������������       �                     $@        e       h                    �?П[;U��?             =@       f       g                 @3�/@���!pc�?             6@        ������������������������       �r�q��?             (@        ������������������������       ����Q��?             $@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KKiKK��h\�B�       �{@      q@     0w@     �V@      @      0@              .@      @      �?     �v@     �R@     �B@      6@       @      @     �A@      1@      3@      @      0@      &@      ,@       @       @      @      (@      @      "@       @      @      @       @      @     �t@     �J@     `o@      >@      X@      6@     �V@      1@     @T@      *@      $@             �Q@      *@      ,@             �L@      *@      K@      @      &@      @      @      @      @             �E@       @       @       @     �A@              @      @      "@      @      @      @      @      �?      @      @     `c@       @      O@      @      M@      @     �F@      @      @@      �?      "@      �?      7@              *@       @      @      �?       @      �?      *@              @       @     @W@      @     @V@       @     �I@       @     �G@      �?      @      �?      C@              @      �?     �S@      7@     �C@      5@      B@      .@      $@      &@      "@      @      �?      @      :@      @      2@      @      $@      �?       @      @       @              @      @     �C@       @      $@       @      =@             @Q@     �f@      B@     �D@              7@      B@      2@              @      B@      (@      0@      $@      @      "@      *@      �?      @      �?      "@              4@       @      @       @      *@             �@@     �a@      0@      9@      1@     �\@      @     �X@      @      =@      �?      9@      �?      $@              .@       @      @      �?     �Q@             �K@      �?      .@      �?      @              $@      *@      0@      @      0@       @      $@      @      @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ� �NhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKuhth)h,K ��h.��R�(KKu��h{�B@         L                    �?�6��l�?�           @�@              7                    �?2�Bo��?(           �{@    @A@                          �:@��h��?�            �t@      5@                           �?���N8�?7             U@       @                            @"pc�
�?	             &@      @������������������������       �      �?             @      @������������������������       �؇���X�?             @      .@       	                   �@��pBI�?.            @R@      @������������������������       �      �?             @      @
                        ���$@@	tbA@�?*            @Q@     �?������������������������       �                     I@     (@                           &@�}�+r��?             3@       @������������������������       �z�G�z�?             @      [@������������������������       �                     ,@      R@       .                 ��$:@d�6��:�?�            @o@     $@       -                 ���+@�׾���?}             h@     @       &                    $@<���D�?m            �d@                               s�@P�R�`M�?X            ``@                               033@ ���J��?            �C@                                 �>@�8��8��?             (@       ������������������������       �z�G�z�?             @n      ������������������������       �                     @�      ������������������������       �                     ;@�                                 �?�A����?<             W@                               ��(@8�Z$���?             :@                                 >@r�q��?             2@      ������������������������       ��q�q�?             "@      ������������������������       �                     "@      ������������������������       �      �?              @�                                �@��IF�E�?,            �P@       ������������������������       �և���X�?             @V              !                   �>@ ,��-�?'            �M@      ������������������������       �                     <@3      "       #                   @@@��� ��?             ?@       ������������������������       ��q�q�?             @�       $       %                   @C@HP�s��?             9@       ������������������������       �                     .@v       ������������������������       �z�G�z�?             $@j       '       (                   �<@������?             A@        ������������������������       �X�<ݚ�?             "@�       )       ,                   @D@�J�4�?             9@       *       +                 `fF)@��S�ۿ?	             .@        ������������������������       �                     @$       ������������������������       �ףp=
�?             $@       ������������������������       ��z�G��?             $@       ������������������������       �                     <@-       /       2                    �?���b���?!            �L@        0       1                 �D8H@R�}e�.�?             :@       ������������������������       �և���X�?             ,@A       ������������������������       ��8��8��?             (@�       3       6                   �I@�g�y��?             ?@       4       5                 `fF<@�q�q�?             5@        ������������������������       �؇���X�?             @�       ������������������������       �և���X�?	             ,@      ������������������������       �z�G�z�?             $@�       8       K                    @������?S            @[@      9       D                     @�lg����?B            �U@      :       ?                    �?Rg��J��?&            �H@      ;       >                     �?��}*_��?             ;@      <       =                   @B@��.k���?             1@       ������������������������       �X�<ݚ�?             "@7      ������������������������       �      �?              @G       ������������������������       �z�G�z�?             $@      @       A                   �:@8�A�0��?             6@       ������������������������       �                     @�      B       C                 `f�R@���Q��?             .@      ������������������������       �      �?              @8       ������������������������       �և���X�?             @8      E       F                    ,@���"͏�?            �B@       ������������������������       �                     @-      G       H                 �&B@��S�ۿ?             >@       ������������������������       �z�G�z�?             @�      I       J                    7@`2U0*��?             9@        ������������������������       �      �?             @�       ������������������������       �                     5@v      ������������������������       �                     7@�      M       l                   �>@f����?�            �p@      N       i                    @�qǩ�?s             h@      O       d                 039@����!��?e             f@      P       W                    �?���b���?C            �\@       Q       V                 ��.@      �?             F@       R       U                   P,@�!���?             A@      S       T                 ��|$@�J�4�?             9@      ������������������������       �������?
             1@%      ������������������������       �                      @g      ������������������������       ��<ݚ�?             "@�       ������������������������       �                     $@y       X       [                     @      �?*            �Q@        Y       Z                   �9@z�G�z�?
             .@        ������������������������       �؇���X�?             @        ������������������������       �      �?              @        \       a                   �;@<|ۤ$�?             �K@       ]       `                    �?��
ц��?            �C@       ^       _                   �7@�q�q�?             8@       ������������������������       ���S���?             .@        ������������������������       ��<ݚ�?             "@        ������������������������       �������?             .@        b       c                 @3#%@      �?
             0@        ������������������������       �                     @        ������������������������       �z�G�z�?             $@        e       h                 03�a@X��Oԣ�?"             O@       f       g                    �? "��u�?             I@       ������������������������       �                     D@        ������������������������       ��z�G��?             $@        ������������������������       ��q�q�?             (@        j       k                   �3@      �?             0@        ������������������������       �                     @        ������������������������       �X�<ݚ�?             "@        m       n                   @C@�S(��d�?5            @S@        ������������������������       �                    �@@        o       t                    @��2(&�?             F@       p       q                   �H@ ���J��?            �C@       ������������������������       �                     :@        r       s                     �?$�q-�?             *@       ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �t�b�      h�h)h,K ��h.��R�(KKuKK��h\�BP       0{@     Pq@     �v@     �S@     �q@     �G@      T@      @      "@       @      @      �?      @      �?     �Q@       @      @      �?      Q@      �?      I@              2@      �?      @      �?      ,@             �i@     �E@     �e@      4@      b@      4@     �]@      (@      C@      �?      &@      �?      @      �?      @              ;@             @T@      &@      6@      @      .@      @      @      @      "@              @      �?     �M@      @      @      @     �K@      @      <@              ;@      @      @       @      7@       @      .@               @       @      :@       @      @      @      5@      @      ,@      �?      @              "@      �?      @      @      <@              A@      7@      3@      @       @      @      &@      �?      .@      0@      @      ,@      �?      @      @       @       @       @     @S@      @@      K@      @@      :@      7@      1@      $@      "@       @      @      @      @      @       @       @      "@      *@              @      "@      @      @       @      @      @      <@      "@              @      <@       @      @      �?      8@      �?      @      �?      5@              7@             �Q@     �h@     @P@     �_@     �J@     �^@      G@      Q@      &@     �@@      &@      7@      @      5@      @      *@               @      @       @              $@     �A@     �A@      @      (@      �?      @       @      @      @@      7@      2@      5@      ,@      $@      @       @      @       @      @      &@      ,@       @      @               @       @      @     �K@      @     �G@              D@      @      @      @       @      (@      @      @              @      @      @     �Q@             �@@      @      C@      �?      C@              :@      �?      (@      �?      @              @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ���bhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKihth)h,K ��h.��R�(KKi��h{�B@         P                    �?\H�l�?�           @�@                                  @�,��h�?6           0~@ �x                              @�d�����?             3@     &@������������������������       �        	             *@        ������������������������       �r�q��?             @      �?                            �?����?(            }@      &@                          �9@�û��|�?9             W@        ������������������������       �                     @      @	                        ��";@�ģ�a@�?4            @U@       @
                          �H@p�ݯ��?	             3@     @������������������������       ��q�q�?             (@      �?������������������������       �և���X�?             @      @                          @B@���|���?+            �P@     ,@                          �@@�s��:��?             C@     @@������������������������       �f���M�?             ?@       @������������������������       �؇���X�?             @      *@                           �?      �?             <@       ������������������������       ����Q��?             $@�                                 �?r�q��?             2@       ������������������������       �                     @w                              03�U@      �?
             (@      ������������������������       �؇���X�?             @�      ������������������������       ����Q��?             @�             O                 �T�I@��r
'��?�            @w@             N                    �?����@��?�            �v@             C                 ���+@�Yr8{�?�            pu@                                  �?�¤�hJ�?�             q@                                 �7@�������?             >@       ������������������������       ����Q��?             @�                                @<@�J�4�?             9@      ������������������������       �������?	             1@V      ������������������������       �                      @J      !       4                   �<@�������?�            @n@      "       3                    �?�C��H�?g            `c@      #       $                   �2@�M�N���?`            @b@        ������������������������       �        
             3@�       %       (                   �3@L<8)��?V            �_@        &       '                 �?�@r�q��?             2@       ������������������������       �                      @�       ������������������������       ��z�G��?             $@�       )       *                    �?��Ujѡ�?K            @[@        ������������������������       �                     1@�       +       ,                 �1@���.�6�?@             W@        ������������������������       �؇���X�?             <@       -       .                 pf� @      �?+             P@       ������������������������       �                    �D@-       /       0                    $@���}<S�?             7@        ������������������������       ������H�?             "@�       1       2                   �:@@4և���?	             ,@       ������������������������       �                     "@�       ������������������������       �z�G�z�?             @�       ������������������������       ��q�q�?             "@�       5       :                 �?�@��{H�?9            �U@        6       7                 ���@ >�֕�?            �A@       ������������������������       �        
             .@�       8       9                    A@ףp=
�?             4@       ������������������������       �"pc�
�?             &@:      ������������������������       �                     "@;      ;       <                 @3�@�θ�?"             J@       ������������������������       ��eP*L��?             &@I      =       >                 ���"@�p ��?            �D@       ������������������������       ���S�ۿ?             .@G       ?       @                   �'@���B���?             :@       ������������������������       ��	j*D�?             *@!      A       B                   @D@$�q-�?             *@       ������������������������       �                     "@�      ������������������������       �      �?             @8       D       G                   �4@0z�(>��?+            �Q@       E       F                 03;4@z�G�z�?             $@       ������������������������       �z�G�z�?             @-      ������������������������       �z�G�z�?             @,      H       I                 039@��v$���?#            �N@      ������������������������       �                     B@�       J       K                    �?`2U0*��?             9@        ������������������������       �                     "@v      L       M                 0C\;@      �?	             0@       ������������������������       �؇���X�?             @�      ������������������������       �                     "@�      ������������������������       �                     3@�      ������������������������       ����Q��?             $@�      Q       d                    �?j[j�v��?�            �l@       R       W                 `fV$@�:�B��?r             f@       S       T                   �9@�e����?            �C@       ������������������������       ��G��l��?             5@%      U       V                    �?�E��ӭ�?             2@       ������������������������       �r�q��?             @�       ������������������������       ��q�q�?             (@y       X       _                   �<@�θV�?Y            @a@        Y       Z                     @z�G�z�?'             N@       ������������������������       �                    �A@        [       \                   �&@�q�����?             9@        ������������������������       �      �?              @        ]       ^                    �?j���� �?             1@        ������������������������       �                     @        ������������������������       ��q�q�?             (@        `       a                   �H@ ���J��?2            �S@       ������������������������       �        &             O@        b       c                    J@      �?             0@        ������������������������       ��q�q�?             @        ������������������������       �                     $@        e       f                 `v�6@$��m��?             J@        ������������������������       �X�Cc�?             ,@        g       h                     @�I�w�"�?             C@        ������������������������       �                      @        ������������������������       �(;L]n�?             >@        �t�bh�h)h,K ��h.��R�(KKiKK��h\�B�       �|@     �o@     �x@     �V@      @      ,@              *@      @      �?     @x@      S@      L@      B@      @             �H@      B@      @      (@      @       @      @      @      E@      8@      5@      1@      4@      &@      �?      @      5@      @      @      @      .@      @      @              "@      @      @      �?      @       @     �t@      D@     `t@      B@     0s@      B@     �m@     �@@      7@      @       @      @      5@      @      *@      @       @              k@      :@     �a@      (@      a@      "@      3@             �]@      "@      .@      @       @              @      @     �Y@      @      1@             �U@      @      8@      @      O@       @     �D@              5@       @       @      �?      *@      �?      "@              @      �?      @      @     @R@      ,@     �@@       @      .@              2@       @      "@       @      "@              D@      (@      @      @     �A@      @      ,@      �?      5@      @      "@      @      (@      �?      "@              @      �?      Q@      @       @       @      @      �?      @      �?      N@      �?      B@              8@      �?      "@              .@      �?      @      �?      "@              3@              @      @      P@     �d@      >@     `b@      0@      7@      &@      $@      @      *@      �?      @      @       @      ,@      _@      (@      H@             �A@      (@      *@       @      @      $@      @      @              @      @       @      S@              O@       @      ,@       @      @              $@      A@      2@      @      "@      =@      "@               @      =@      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ+�MhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKahth)h,K ��h.��R�(KKa��h{�B@         $                 �=/@�JX-��?�           @�@                               `f�$@�[%�r�?�            �w@      �                           �?؇���X�?�            q@                                  �7@�E��ӭ�?/             R@      �?                          �4@��S���?	             .@     6@������������������������       �      �?             @      *@������������������������       �X�<ݚ�?             "@      @                          @<@���y4F�?&            �L@      @	                           �?���!pc�?             F@     @
                           �? 7���B�?             ;@      @������������������������       �                     $@      �?������������������������       ��IєX�?             1@      �?������������������������       �ҳ�wY;�?
             1@       @������������������������       �                     *@                                   �?�j�zZ��?�             i@     .@                          �8@�IєX�?r            @e@      @                          �0@p���?#             I@       ������������������������       �r�q��?             @�      ������������������������       �                     F@�                                  @��(\���?O             ^@       ������������������������       �                     *@n                              ��@ܑ-Z���?H            �Z@       ������������������������       ����Q��?             @�      ������������������������       ��v�\�?D            �Y@�                              @3�@¦	^_�?             ?@                               �&B@��S���?             .@       ������������������������       �X�<ݚ�?             "@      ������������������������       ��q�q�?             @      ������������������������       �      �?             0@�                              ���+@xZ�l ��??            �Z@      ������������������������       ����=�/�?)            @Q@V              !                    �?�˹�m��?             C@      ������������������������       �                     6@3      "       #                    �?     ��?
             0@      ������������������������       �      �?              @�       ������������������������       �      �?              @�       %       N                    �?����n��?�            �t@       &       )                 ��`3@Ks��?p            �f@        '       (                    �?X�<ݚ�?	             2@       ������������������������       ������H�?             "@�       ������������������������       �                     "@�       *       -                 03�9@�4�t���?g            `d@        +       ,                    �? �q�q�?             8@       ������������������������       �        	             1@       ������������������������       �؇���X�?             @       .       K                    @�x��j��?Y            `a@       /       0                    #@�5C�z�?H            �\@        ������������������������       �                     @�       1       B                   @C@�Sb(�	�?D             [@       2       ;                    �?j���� �?(             Q@       3       6                   �>@��Q��?             D@        4       5                 03k:@�eP*L��?             &@        ������������������������       �      �?             @�       ������������������������       �����X�?             @      7       :                    >@�c�Α�?             =@       8       9                   `F@ףp=
�?             4@       ������������������������       �؇���X�?             @:      ������������������������       �$�q-�?             *@;      ������������������������       ��q�q�?             "@?      <       ?                     �?      �?             <@       =       >                    �?������?             .@       ������������������������       �      �?              @G       ������������������������       �؇���X�?             @      @       A                 0C�:@�θ�?             *@       ������������������������       �      �?              @�      ������������������������       �                     @�      C       H                 03�>@z�G�z�?             D@        D       G                     �?���!pc�?             6@      E       F                 `f�;@ҳ�wY;�?	             1@      ������������������������       ��<ݚ�?             "@-      ������������������������       �      �?              @,      ������������������������       �                     @�      I       J                    �?�X�<ݺ?             2@        ������������������������       �      �?             @�       ������������������������       �                     ,@v      L       M                 ���A@`2U0*��?             9@       ������������������������       �r�q��?             @�      ������������������������       �                     3@�      O       Z                    �?.�*���?_            �b@      P       Y                    @�S#א��?E            @]@      Q       X                 03[=@�8��8��?A             [@        R       S                    :@�θ�?            �C@       ������������������������       �        
             2@-      T       U                   �>@և���X�?             5@       ������������������������       �      �?              @g      V       W                   @G@�	j*D�?	             *@       ������������������������       �                     @y       ������������������������       �      �?              @}       ������������������������       �        *            @Q@�       ������������������������       �X�<ݚ�?             "@        [       `                    ?@      �?             A@       \       ]                    �?���Q��?             9@        ������������������������       ��z�G��?             $@        ^       _                    @z�G�z�?             .@        ������������������������       ����Q��?             @        ������������������������       �ףp=
�?             $@        ������������������������       ��<ݚ�?             "@        �t�bh�h)h,K ��h.��R�(KKaKK��h\�B       @}@     �n@     Ps@     �Q@     @m@     �C@      J@      4@      @       @      @      @      @      @     �F@      (@      @@      (@      :@      �?      $@              0@      �?      @      &@      *@             �f@      3@      d@      $@     �H@      �?      @      �?      F@             �[@      "@      *@             �X@      "@      @       @     �W@      @      6@      "@       @      @      @      @      @       @      ,@       @     �R@      @@      D@      =@     �A@      @      6@              *@      @      @       @      @      �?     �c@     �e@      `@     �J@       @      $@       @      �?              "@      ^@     �E@      7@      �?      1@              @      �?     @X@      E@     @R@     �D@              @     @R@     �A@      D@      <@      :@      ,@      @      @      @      �?       @      @      5@       @      2@       @      @      �?      (@      �?      @      @      ,@      ,@      @      &@      @      @      �?      @      $@      @      @      @      @             �@@      @      0@      @      &@      @      @       @      @      @      @              1@      �?      @      �?      ,@              8@      �?      @      �?      3@              ?@      ^@      ,@     �Y@      "@     �X@      "@      >@              2@      "@      (@      @      @      @      "@              @      @      @             @Q@      @      @      1@      1@      .@      $@      @      @      (@      @      @       @      "@      �?       @      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJY]hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKkhth)h,K ��h.��R�(KKk��h{�B�         N                    �?��!h
��?�           @�@              3                 ��i=@�q�q�?5            ~@              2                    @R�f?���?�            @w@     @@                           !@��Ns��?�            �v@      �?������������������������       �                      @     6@                          �;@d{̯E>�?�            `v@      *@                          �:@J3�xH��?N             `@     @       	                 ���@�(�,�J�?I            �]@       @������������������������       ��eP*L��?             &@     @
                          �5@ ˤ���?A            �Z@     @                        ��Y @����|e�?%             K@     �?                        �?�@:ɨ��?            �@@     �?                        �1@�q�q�?             8@      @                         s�@�q�q�?	             .@       ������������������������       �؇���X�?             @     .@������������������������       �      �?              @      @������������������������       �                     "@Z      ������������������������       �X�<ݚ�?             "@�                              ���$@؇���X�?             5@       ������������������������       �                     $@w                                  @���!pc�?	             &@       ������������������������       �z�G�z�?             @�      ������������������������       ��q�q�?             @�                                �8@�O4R���?            �J@      ������������������������       �                     A@�                              �?�@�}�+r��?             3@       ������������������������       �r�q��?             @      ������������������������       �                     *@      ������������������������       ����|���?             &@�             !                     �?��F!�?�            �l@                                ��$:@�>4և��?             <@       ������������������������       �                     "@J      ������������������������       ��d�����?             3@3      "       1                   @E@�qM�R��?�             i@      #       $                 �?�@xif�N��?o            �e@        ������������������������       �Х-��ٹ?4            �R@�       %       &                 @3�@؇���X�?;            �X@        ������������������������       ��q�q�?             (@j       '       ,                 `��+@���W���?5            �U@        (       )                     @z�G�z�?             D@        ������������������������       �X�<ݚ�?             "@�       *       +                   �=@��a�n`�?             ?@        ������������������������       �d}h���?	             ,@$       ������������������������       �        	             1@       -       .                    �?�nkK�?             G@        ������������������������       �        
             2@-       /       0                   �<@@4և���?             <@        ������������������������       ��<ݚ�?             "@�       ������������������������       �                     3@A       ������������������������       �                     <@�       ������������������������       �                     @�       4       7                    !@���B��?G             [@        5       6                 �D C@����X�?             ,@        ������������������������       �      �?              @      ������������������������       �      �?             @�       8       9                    /@6n�
$)�??            �W@       ������������������������       �                     "@:      :       I                    �?Ї?��f�?:            @U@      ;       H                     @���>4��?'             L@      <       G                     �?�q�q��?#             H@      =       B                 �!�I@D^��#��?            �D@      >       ?                    �?�q�q�?             ;@        ������������������������       �      �?             $@      @       A                   �<@������?             1@      ������������������������       ��z�G��?             $@�      ������������������������       �؇���X�?             @�      C       D                    >@����X�?             ,@        ������������������������       ����Q��?             @8      E       F                   @G@�<ݚ�?             "@       ������������������������       �z�G�z�?             @-      ������������������������       �      �?             @,      ������������������������       �                     @�      ������������������������       �      �?              @�       J       K                 ���S@>���Rp�?             =@       ������������������������       �        
             *@v      L       M                 `fa@     ��?	             0@      ������������������������       ��q�q�?             "@�      ������������������������       �؇���X�?             @�      O       X                     @>��C��?�             m@      P       S                    6@��*����?U            `a@       Q       R                    �?�L���?            �B@        ������������������������       �                      @      ������������������������       �ܷ��?��?             =@-      T       U                    �?�K}��?>            �Y@       ������������������������       �                     D@g      V       W                 03�a@0�z��?�?(             O@       ������������������������       �        "            �J@y       ������������������������       ������H�?             "@}       Y       h                 ��Y7@ܐ҆��?C            @W@       Z       ]                    �?���Q��?5            �R@        [       \                    �?����>�?            �B@       ������������������������       �z�G�z�?             9@        ������������������������       ��q�q�?             (@        ^       c                    �?�\��N��?             C@       _       `                   �6@r�q��?             8@        ������������������������       ��<ݚ�?             "@        a       b                 ��� @���Q��?             .@       ������������������������       ��<ݚ�?             "@        ������������������������       ��q�q�?             @        d       g                    �?X�Cc�?             ,@       e       f                 ���.@�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       ����Q��?             @        i       j                    @�����H�?             2@        ������������������������       ����Q��?             @        ������������������������       �        
             *@        �t�bh�h)h,K ��h.��R�(KKkKK��h\�B�       �z@     �q@     �w@      Y@     �s@     �L@     Ps@     �L@               @     Ps@     �H@     �Y@      :@     �X@      3@      @      @     @W@      ,@     �D@      *@      7@      $@      3@      @      $@      @      @      �?      @      @      "@              @      @      2@      @      $@               @      @      @      �?      @       @      J@      �?      A@              2@      �?      @      �?      *@              @      @     �i@      7@      7@      @      "@              ,@      @     �f@      2@     `c@      2@     �Q@      @      U@      ,@      @      @     @S@      "@     �@@      @      @      @      <@      @      &@      @      1@              F@       @      2@              :@       @      @       @      3@              <@              @             @P@     �E@      @      $@      �?      @      @      @     �N@     �@@      "@              J@     �@@      >@      :@      =@      3@      6@      3@      2@      "@      @      @      *@      @      @      @      @      �?      @      $@       @      @       @      @      �?      @      �?      @      @              �?      @      6@      @      *@              "@      @      @      @      @      �?      I@     �f@      @     �`@      @      A@               @      @      :@      �?     @Y@              D@      �?     �N@             �J@      �?       @      G@     �G@      >@     �F@      $@      ;@      @      4@      @      @      4@      2@      &@      *@       @      @      "@      @      @       @       @      @      "@      @      @       @      @               @       @       @      @      0@       @      @       @      *@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ4
hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKghth)h,K ��h.��R�(KKg��h{�B�         H                    �?������?�           @�@                                  �?�Sn��?*           �}@  ute th                          @@j����?9            �T@                                ���@�����H�?             2@ �>	�  ������������������������       �                      @     6@������������������������       �z�G�z�?             $@      *@                           4@���Q��?)            @P@      @������������������������       �      �?              @       @	                         I>@p�ݯ��?%            �L@      @
                        @Q,@�+e�X�?             9@      @������������������������       �և���X�?             @     �?������������������������       ������H�?             2@     �?                        @�pX@     ��?             @@      @                        pVAH@b�2�tk�?             2@        ������������������������       �      �?              @     .@������������������������       ��z�G��?             $@      @                           �?����X�?             ,@       ������������������������       ��z�G��?             $@�      ������������������������       �      �?             @�                                  �?��|��?�            `x@                               03�U@����0�?#             K@                                �J@���!pc�?             F@                              ���M@ҳ�wY;�?             A@                                �9@X�<ݚ�?             ;@       ������������������������       �                     @�      ������������������������       ��eP*L��?             6@c      ������������������������       �                     @      ������������������������       �                     $@      ������������������������       ��z�G��?             $@�             -                 @3�@ �Cc}�?�             u@              ,                   @F@�?�'�@�?\             c@              )                 �?�@��ED���?R             `@      !       "                   �7@X�
����?I             ]@       ������������������������       �������?             B@A      #       (                 �{@z�G�z�?5             T@       $       '                    �?�������?'             N@        %       &                   �<@ףp=
�?             4@       ������������������������       ���S�ۿ?
             .@j       ������������������������       �z�G�z�?             @�       ������������������������       ��z�G��?             D@�       ������������������������       �                     4@�       *       +                   �?@�n_Y�K�?	             *@        ������������������������       �      �?             @$       ������������������������       �����X�?             @       ������������������������       �        
             7@       .       A                    �?���}<S�?r             g@       /       0                    �?�5[|/��?R            �`@        ������������������������       �؇���X�?             @�       1       6                    ?@H�Swe�?M            @_@       2       5                 ���!@`׀�:M�?-            �R@        3       4                   �;@      �?             0@        ������������������������       �      �?              @�       ������������������������       �                      @�       ������������������������       �        !             M@      7       @                    �?`�H�/��?             �I@       8       =                     @X�EQ]N�?            �E@      9       :                   �B@�J�4�?             9@       ������������������������       �      �?              @;      ;       <                   @F@�IєX�?             1@       ������������������������       �r�q��?             @I      ������������������������       �                     &@7      >       ?                   �@@�X�<ݺ?             2@        ������������������������       �r�q��?             @      ������������������������       �                     (@!      ������������������������       �                      @�      B       G                    !@D>�Q�?              J@       C       D                     @և���X�?             5@        ������������������������       �                     @8      E       F                 033>@      �?
             0@       ������������������������       ����Q��?             $@-      ������������������������       �                     @,      ������������������������       �                     ?@�      I       N                     @��1+�?�            �m@        J       K                   �H@�Ru߬Α?L            �\@       ������������������������       �        B            @Y@v      L       M                 03[;@$�q-�?
             *@       ������������������������       �                     @�      ������������������������       �؇���X�?             @�      O       V                    �?l��TO��?L            @_@       P       U                 ��.@      �?             J@      Q       R                    �?�q�q�?            �C@        ������������������������       ����Q��?             @      S       T                   �5@�t����?             A@       ������������������������       ��q�q�?             "@%      ������������������������       � �o_��?             9@g      ������������������������       �        	             *@�       W       d                    �?��T���?/            @R@       X       c                   �A@�F�j��?#            �J@       Y       \                   �4@�&!��?            �E@        Z       [                    (@�eP*L��?             &@        ������������������������       ����Q��?             @        ������������������������       ��q�q�?             @        ]       b                    �?     ��?             @@       ^       a                   �;@��+7��?             7@       _       `                    9@r�q��?             2@       ������������������������       �      �?             (@        ������������������������       �                     @        ������������������������       ����Q��?             @        ������������������������       �X�<ݚ�?             "@        ������������������������       �                     $@        e       f                 ��T?@P���Q�?             4@       ������������������������       �                     *@        ������������������������       �؇���X�?             @        �t�bh�h)h,K ��h.��R�(KKgKK��h\�Bp        |@     `p@     `x@     �T@     �K@      <@      0@       @       @               @       @     �C@      :@      @      @      B@      5@      3@      @      @      @      0@       @      1@      .@      @      &@      @      @      @      @      $@      @      @      @      @      �?     �t@     �K@     �A@      3@      @@      (@      6@      (@      .@      (@      @              $@      (@      @              $@              @      @     �r@      B@     �`@      4@     @[@      4@     @Y@      .@     �A@      �?     �P@      ,@      G@      ,@      2@       @      ,@      �?      @      �?      <@      (@      4@               @      @      @      @      @       @      7@              e@      0@     @_@      @      @      �?     �]@      @     @R@      �?      .@      �?      @      �?       @              M@              G@      @      C@      @      5@      @      @      @      0@      �?      @      �?      &@              1@      �?      @      �?      (@               @             �E@      "@      (@      "@              @      (@      @      @      @      @              ?@              N@     `f@      �?     @\@             @Y@      �?      (@              @      �?      @     �M@     �P@      *@     �C@      *@      :@      @       @      $@      8@      @      @      @      2@              *@      G@      ;@      ;@      :@      1@      :@      @      @       @      @      @       @      &@      5@      @      1@      @      .@      @      "@              @      @       @      @      @      $@              3@      �?      *@              @      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��;hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKahth)h,K ��h.��R�(KKa��h{�B@         N                 0�&H@\H�l�?�           @�@                               `f�$@�#�����?d           P�@      @                          �1@
�GN��?�            �p@        ������������������������       ��eP*L��?             6@       @                           �?*��
�?�            @n@     6@                          �;@H"Б$�?y            �h@      *@                           �?� y���?'            �P@     @                        pf� @�r����?#             N@      @	       
                 03�@ףp=
�?             I@      @������������������������       �d}h���?             ,@      @                        @3�@�X�<ݺ?             B@     �?������������������������       �                     4@     �?                          �4@      �?             0@       @������������������������       �"pc�
�?             &@        ������������������������       �                     @     .@������������������������       ��z�G��?             $@      @������������������������       �և���X�?             @Z                              ���@t��ճC�?R            �`@       ������������������������       �                     A@�                              ���@�)���Y�??            �X@       ������������������������       ��z�G��?             $@n                              pFt @t��ճC�?:             V@      ������������������������       ��S(��d�?3            @S@�      ������������������������       �                     &@�                                �9@X��ʑ��?            �E@                               ���@�q�q�?
             2@       ������������������������       �      �?              @      ������������������������       �ףp=
�?             $@      ������������������������       ����Q��?             9@�             ;                    �?<�m�7�?�             t@             $                    $@Ժe�R�?t            �h@               !                    @      �?             @@      ������������������������       �                     3@3      "       #                    @$�q-�?	             *@       ������������������������       �r�q��?             @�       ������������������������       �                     @�       %       *                     �?�)x��?_            �d@        &       )                   �>@<ݚ)�?             B@       '       (                 �ܵ<@���Q��?             9@       ������������������������       �     ��?             0@�       ������������������������       ��<ݚ�?             "@�       ������������������������       ��C��2(�?             &@�       +       .                    �?x�]AgȽ?I             `@        ,       -                   �<@��s����?             5@       ������������������������       �����X�?             ,@       ������������������������       �                     @-       /       :                    �? 7���B�?=             [@       0       9                   �I@HP�s��?              I@       1       8                     @������?            �D@       2       7                   �*@      �?             @@       3       4                   �;@�8��8��?             8@        ������������������������       �                     $@�       5       6                    @@؇���X�?
             ,@        ������������������������       ��q�q�?             @      ������������������������       �                      @�       ������������������������       �                      @`      ������������������������       �                     "@:      ������������������������       ��<ݚ�?             "@;      ������������������������       �                     M@?      <       A                     @���k�6�?U            @_@      =       @                    6@P���Q�?,             N@       >       ?                   `1@ �Cc}�?             <@       ������������������������       �                     5@      ������������������������       �և���X�?             @!      ������������������������       �                     @@�      B       K                    �?�G\�c�?)            @P@      C       J                 ���4@�Gi����?            �B@       D       G                   �:@����X�?             <@       E       F                 ���,@�eP*L��?             &@       ������������������������       �      �?             @-      ������������������������       �և���X�?             @,      H       I                 ��Y/@�t����?             1@      ������������������������       ��<ݚ�?             "@�       ������������������������       �                      @�       ������������������������       ��<ݚ�?             "@v      L       M                    �?�>4և��?             <@       ������������������������       �      �?             $@�      ������������������������       �        
             2@�      O       ^                    �?X�Cc�?Q            �_@       P       S                   �;@���h%��?(            �O@       Q       R                    �?X�Cc�?	             ,@       ������������������������       �      �?              @      ������������������������       ��q�q�?             @-      T       W                    �?���c�H�?            �H@       U       V                 @�pX@��Q��?             4@      ������������������������       �X�<ݚ�?             "@�       ������������������������       �"pc�
�?             &@y       X       ]                 `fJT@\-��p�?             =@       Y       \                    �?���}<S�?             7@       Z       [                   �@@�r����?
             .@       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       ��q�q�?             @        _       `                    �?�i�y�?)            �O@       ������������������������       �        !            �I@        ������������������������       �r�q��?             (@        �t�bh�h)h,K ��h.��R�(KKaKK��h\�B       �|@     �o@     �y@     �e@     �j@     �I@      (@      $@      i@     �D@     `f@      4@      L@      &@      J@       @     �F@      @      &@      @      A@       @      4@              ,@       @      "@       @      @              @      @      @      @     �^@      "@      A@             @V@      "@      @      @     �T@      @     �Q@      @      &@              6@      5@      (@      @      @      @      "@      �?      $@      .@     �h@     �^@     �c@     �C@      (@      4@              3@      (@      �?      @      �?      @             @b@      3@      9@      &@      .@      $@      *@      @       @      @      $@      �?     @^@       @      1@      @      $@      @      @              Z@      @      G@      @     �C@       @      >@       @      6@       @      $@              (@       @      @       @       @               @              "@              @       @      M@             �D@      U@      @     �L@      @      9@              5@      @      @              @@      C@      ;@      .@      6@       @      4@      @      @       @       @      @      @       @      .@       @      @               @      @       @      7@      @      @      @      2@             �F@     @T@     �E@      4@      @      "@      �?      @      @       @      C@      &@      *@      @      @      @      "@       @      9@      @      5@       @      *@       @      @       @      @               @              @       @       @     �N@             �I@       @      $@�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJS�)/hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsK�hth)h,K ��h.��R�(KK���h{�B�          r                 03�I@�1�uџ�?�           @�@              O                    �?<Z���?{           X�@      @       B                    �?P�b����?           0z@     �?       ;                 ��=@4�|F�?�            �v@      @                           �?��E�B��?�            �t@      6@                        м;4@��[�p�?            �G@     *@       
                   �=@      �?             D@     @       	                    ;@�4�����?             ?@       @������������������������       ��eP*L��?             &@      @������������������������       �      �?             4@      @������������������������       �                     "@     �?������������������������       �                     @     �?       2                    �?Tri����?�            �q@      @                         ��@�����H�?�            `n@                                ���@`���i��?             F@      .@������������������������       �                     7@      @                        ���@���N8�?             5@       ������������������������       �      �?             @�      ������������������������       �        
             1@�                                  �?���\��?�            �h@                                  H@8�Z$���?	             *@      ������������������������       �      �?              @�      ������������������������       �z�G�z�?             @�             1                   �*@��� ��?|            @g@                                �3@Р�31�?q             e@                                 �2@������?             >@                                �0@r�q��?             8@       ������������������������       ��q�q�?             (@      ������������������������       �                     (@�      ������������������������       ��q�q�?             @(             "                     @dҁ
_�?`            `a@               !                   �@@؇���X�?             5@       ������������������������       �                     &@3      ������������������������       ��z�G��?             $@A      #       ,                   �>@�!���?P            �]@       $       %                    �?�c:��?8             W@        ������������������������       �8�Z$���?             *@v       &       '                   �:@86��Z�?0            �S@        ������������������������       �                     =@�       (       +                   �<@ףp=
�?             I@       )       *                 ��) @�Ra����?             F@       ������������������������       ��˹�m��?             C@�       ������������������������       ��q�q�?             @$       ������������������������       �                     @       -       .                   @@@�θ�?             :@        ������������������������       �      �?              @-       /       0                   @C@�����H�?             2@        ������������������������       �                     @�       ������������������������       �"pc�
�?
             &@A       ������������������������       �                     1@�       3       4                    �?�ݜ�?            �C@        ������������������������       ����!pc�?             &@�       5       :                   �@@@4և���?             <@       6       7                     @ףp=
�?             4@       ������������������������       �      �?             @�       8       9                   �:@      �?
             0@       ������������������������       �r�q��?             @:      ������������������������       �                     $@;      ������������������������       �                      @?      <       A                 `f�B@�E��ӭ�?             B@      =       >                    @@���Q��?             9@       ������������������������       �X�<ݚ�?             "@G       ?       @                   �K@     ��?	             0@      ������������������������       �؇���X�?             @!      ������������������������       �X�<ݚ�?             "@�      ������������������������       �                     &@�      C       F                     @����|e�?&             K@        D       E                    /@��
ц��?
             *@       ������������������������       �                     @      ������������������������       �                     @-      G       L                    �?�p ��?            �D@      H       I                    @ �Cc}�?             <@       ������������������������       ��<ݚ�?             "@�       J       K                    3@�}�+r��?             3@        ������������������������       �                     "@v      ������������������������       �ףp=
�?             $@�      M       N                    @�θ�?
             *@       ������������������������       �      �?             @�      ������������������������       �                     @�      P       ]                 `f�$@,Tg�x��?j             e@       Q       R                 ���@�n_Y�K�?"             J@        ������������������������       �      �?             (@      S       V                   �5@��Q���?             D@       T       U                 @� @��S�ۿ?             .@       ������������������������       �      �?              @g      ������������������������       �                     @�       W       X                 �̌@���Q��?             9@        ������������������������       �X�<ݚ�?             "@}       Y       \                   �<@     ��?             0@       Z       [                    ;@"pc�
�?             &@        ������������������������       �����X�?             @        ������������������������       �                     @        ������������������������       ����Q��?             @        ^       g                    �?�������?H             ]@       _       b                 P�>,@     8�?'             P@       `       a                   �9@�C��2(�?            �@@        ������������������������       ����!pc�?             &@        ������������������������       �                     6@        c       d                 ��80@r֛w���?             ?@        ������������������������       �r�q��?             @        e       f                 03�7@H%u��?             9@        ������������������������       �                     $@        ������������������������       �z�G�z�?             .@        h       i                    �?��
ц��?!             J@        ������������������������       �d}h���?
             ,@        j       m                   �9@�s��:��?             C@        k       l                    �?�n_Y�K�?	             *@        ������������������������       �                     @        ������������������������       �r�q��?             @        n       q                    �?��H�}�?             9@       o       p                 0339@      �?
             4@        ������������������������       �                     &@        ������������������������       �X�<ݚ�?             "@        ������������������������       �z�G�z�?             @        s       |                    �?2]��a�?N            @_@        t       {                     @��WV��?              J@       u       v                    �?��
ц��?            �C@        ������������������������       ���
ц��?             *@        w       x                 03�M@
j*D>�?             :@        ������������������������       ������H�?             "@        y       z                    �?j���� �?             1@        ������������������������       �      �?              @        ������������������������       ��<ݚ�?             "@        ������������������������       ��n_Y�K�?             *@        }       ~                    �?0�й���?.            @R@       ������������������������       �        !            �I@               �                 ���W@8�A�0��?             6@        ������������������������       �      �?              @        �       �                 Ъ�c@d}h���?             ,@        ������������������������       �      �?              @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��h\�B0       P|@     0p@     Pz@     �d@      v@     @P@     �s@      J@     �q@      E@     �B@      $@      >@      $@      5@      $@      @      @      .@      @      "@              @             @o@      @@      k@      ;@     �E@      �?      7@              4@      �?      @      �?      1@             �e@      :@      &@       @      @      �?      @      �?     @d@      8@      b@      8@      6@       @      4@      @       @      @      (@               @      @     �^@      0@      2@      @      &@              @      @     @Z@      *@     @U@      @      &@       @     �R@      @      =@             �F@      @     �C@      @     �A@      @      @       @      @              4@      @      @      @      0@       @      @              "@       @      1@              A@      @       @      @      :@       @      2@       @      @      �?      .@      �?      @      �?      $@               @              :@      $@      .@      $@      @      @      &@      @      @      �?      @      @      &@             �D@      *@      @      @              @      @             �A@      @      9@      @      @       @      2@      �?      "@              "@      �?      $@      @      @      @      @             �P@     @Y@      @@      4@      @      "@      =@      &@      ,@      �?      @      �?      @              .@      $@      @      @      &@      @      "@       @      @       @      @               @      @     �A@     @T@      &@     �J@      @      >@      @       @              6@       @      7@      @      �?      @      6@              $@      @      (@      8@      <@      @      &@      5@      1@      @       @              @      @      �?      0@      "@      .@      @      &@              @      @      �?      @      @@     @W@      7@      =@      2@      5@      @      @      &@      .@      �?       @      $@      @      @      @      @       @      @       @      "@      P@             �I@      "@      *@      @       @      @      &@      @      @              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ[س=hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKqhth)h,K ��h.��R�(KKq��h{�B@         N                    �?l��n�?�           @�@              '                 ��l1@��.D��?0           P~@     $@                        �?�@��
CJ�?�            `r@      *@                          �=@ףp=
�?Z            �b@     @       
                   �7@������?C             \@      6@                          �4@      �?             @@     *@������������������������       �        
             3@     @       	                 @�@$�q-�?	             *@      @������������������������       �                      @      @������������������������       �z�G�z�?             @      @                          �;@z�G�z�?0             T@      �?������������������������       �j���� �?             1@     �?                         s�@�����H�?%            �O@       @������������������������       �                     :@                                �?$@��G���?            �B@      .@������������������������       ����Q��?
             .@      @                           �?���7�?             6@        ������������������������       �؇���X�?             @        ������������������������       �                     .@      @������������������������       �                     C@      �?                        @3�@<ݚ��?`             b@      $@������������������������       �      �?             $@      �?                           &@�Y����?Z            �`@      @������������������������       �                     @      @                          �3@��7PB��?U            �_@      �?                          �2@���|���?	             &@    @Y@������������������������       �z�G�z�?             @      �?������������������������       �      �?             @      @                           $@��Õty�?L             ]@        ������������������������       �D>�Q�?"             J@      >@       &                    �?      �?*             P@     �?        !                    �?P���Q�?&             N@      <@������������������������       �r�q��?             @3      "       %                    �? 7���B�?"             K@      #       $                   @D@���N8�?             E@       ������������������������       �Pa�	�?            �@@�       ������������������������       ������H�?             "@v       ������������������������       �                     (@j       ������������������������       �      �?             @�       (       A                  x#J@�ߎx���?v            �g@       )       @                   �C@l��э�?R            �_@       *       ?                 �TaA@X�Cc�?C            �X@       +       2                     �?P*L�9�?<             V@        ,       -                    �?և���X�?            �A@        ������������������������       �r�q��?             @       .       1                 `f�;@l��[B��?             =@       /       0                   �E@b�2�tk�?
             2@        ������������������������       �      �?             @�       ������������������������       ��q�q�?             (@A       ������������������������       ����!pc�?             &@�       3       <                    :@�T`�[k�?&            �J@       4       5                    �?:ɨ��?            �@@        ������������������������       �      �?             @�       6       9                    �?������?             ;@      7       8                 039@$�q-�?             *@       ������������������������       �                     "@`      ������������������������       �      �?             @:      :       ;                 �̜6@և���X�?
             ,@      ������������������������       �      �?              @?      ������������������������       �      �?             @I      =       >                  �=@ףp=
�?             4@      ������������������������       �                     ,@G       ������������������������       ��q�q�?             @      ������������������������       �z�G�z�?             $@!      ������������������������       �                     =@      �?B       M                     @     ��?$             P@     �?C       D                 p��K@����0�?              K@      �?������������������������       �      �?              @      �?E       L                    �?��+7��?             G@     �?F       I                   �B@�θ�?            �C@      �?G       H                   �=@�q�q�?
             (@     �?������������������������       �؇���X�?             @      �?������������������������       �z�G�z�?             @      �?J       K                    �?PN��T'�?             ;@      �?������������������������       ��z�G��?             $@      �?������������������������       ��IєX�?             1@      �?������������������������       �և���X�?             @      �?������������������������       ��z�G��?             $@      �?O       n                    @��'�e��?�            `l@     �?P       i                    �?*��B��?�            �j@     �?Q       `                   �;@������?v            �f@      �?R       ]                    �?�t����?*             Q@     �?S       X                     @�q�q��?             H@      �?T       U                   �7@�θ�?             :@      �?������������������������       �                      @      �?V       W                 ��m1@�q�q�?             2@      �?������������������������       �X�<ݚ�?             "@      �?������������������������       ��<ݚ�?             "@      �?Y       Z                 �&B@8�A�0��?             6@      �?������������������������       �      �?              @        [       \                    5@X�Cc�?	             ,@       ������������������������       �      �?              @        ������������������������       �      �?             @        ^       _                 �F�)@P���Q�?             4@        ������������������������       �z�G�z�?             @        ������������������������       �                     .@        a       f                     @x�}b~|�?L            �\@       b       c                   �H@`׀�:M�?0            �R@       ������������������������       �        $             N@        d       e                   �J@@4և���?             ,@        ������������������������       �      �?             @        ������������������������       �                     $@        g       h                   �@@R���Q�?             D@       ������������������������       �r�q��?             B@        ������������������������       �      �?             @       j       k                 ��97@*;L]n�?             >@        ������������������������       ��8��8��?             (@        l       m                     @�q�q�?             2@       ������������������������       ����Q��?             $@       ������������������������       �                      @        o       p                    :@�q�q�?	             .@       ������������������������       �և���X�?             @        ������������������������       �      �?              @        �t�bh�h)h,K ��h.��R�(KKqKK��h\�B       {@     pq@     �w@     @Z@     @o@      F@     �`@      .@     @X@      .@      ?@      �?      3@              (@      �?       @              @      �?     �P@      ,@      $@      @      L@      @      :@              >@      @      "@      @      5@      �?      @      �?      .@              C@             �\@      =@      @      @     �[@      8@              @     �[@      1@      @      @      @      �?      @      @     �Y@      *@     �E@      "@      N@      @     �L@      @      @      �?      J@       @      D@       @      @@      �?       @      �?      (@              @      �?     @`@     �N@      W@     �A@     �O@     �A@     �N@      ;@      4@      .@      @      �?      .@      ,@      @      &@      @      @      @       @       @      @     �D@      (@      7@      $@      @      @      4@      @      (@      �?      "@              @      �?       @      @      @      @      @      @      2@       @      ,@              @       @       @       @      =@              C@      :@     �A@      3@      �?      @      A@      (@      >@      "@      @      @      @      �?      �?      @      7@      @      @      @      0@      �?      @      @      @      @     �J@     �e@     �E@      e@      >@      c@      4@      H@      3@      =@      @      4@               @      @      (@      @      @       @      @      *@      "@      @      @      "@      @      @       @      @      @      �?      3@      �?      @              .@      $@      Z@      �?     @R@              N@      �?      *@      �?      @              $@      "@      ?@      @      >@      @      �?      *@      1@      �?      &@      (@      @      @      @       @              $@      @      @      @      @       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJnխphG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKShth)h,K ��h.��R�(KKS��h{�B�         2                    �?z��Y�)�?�           @�@                                  @X���?�?2           �~@     @A@                        @3�4@z�G�z�?             4@      5@������������������������       �                     $@       @                           @���Q��?
             $@      "@������������������������       �                     @      @������������������������       �z�G�z�?             @      @       %                   �C@vsSj��?!           �}@     @	       "                 �U�R@ �/gB�?�            `w@     @
                        ��D:@d��o�t�?�            @v@     @                          �2@��8���?�            �q@      �?������������������������       �                     0@     �?                            �?PN��T'�?�            �p@       @������������������������       �                     (@                                   �?��ED���?�             p@      .@                          @@      �?             <@     @������������������������       ����y4F�?             3@Z      ������������������������       ��q�q�?             "@�                                 �?����u�?�            �l@                                s�@ܷ��?��?             =@       ������������������������       �                      @n                                @'@؇���X�?             5@      ������������������������       �؇���X�?	             ,@�      ������������������������       �؇���X�?             @�      ������������������������       �D|U��@�?x             i@�                                 �?��R[s�?+            �Q@                                �?@�L�lRT�?            �F@      ������������������������       �      �?             B@      ������������������������       ��<ݚ�?             "@�             !                   �;@HP�s��?             9@                                @�F@r�q��?	             (@      ������������������������       �                      @J      ������������������������       �      �?             @3      ������������������������       �        	             *@A      #       $                    �?b�2�tk�?             2@        ������������������������       �      �?              @�       ������������������������       ����Q��?             $@v       &       )                    �?P���Q�?9             Y@        '       (                 �D8H@r�q��?	             (@        ������������������������       �z�G�z�?             @�       ������������������������       �؇���X�?             @�       *       1                    �?�zvܰ?0             V@       +       0                    �?(�5�f��?*            �S@       ,       -                 `fF:@��ɉ�?#            @P@       ������������������������       �                    �J@       .       /                   �L@r�q��?             (@        ������������������������       ��q�q�?             @]       ������������������������       �                     @�       ������������������������       �@4և���?             ,@A       ������������������������       �                     "@�       3       <                     @~�1u���?�            @k@       4       9                  "�b@�7��?J            @]@       5       8                   �;@г�wY;�??            �Y@        6       7                    6@Du9iH��?            �E@       ������������������������       �և���X�?             @�       ������������������������       �                     B@`      ������������������������       �        &            �M@:      :       ;                    �?z�G�z�?             .@      ������������������������       �                     $@?      ������������������������       ����Q��?             @I      =       P                 ���4@h0�����?B            @Y@      >       E                 pF @�n_Y�K�?3            �S@        ?       B                   �7@r٣����?            �@@       @       A                    �?�r����?
             .@      ������������������������       �ףp=
�?             $@      �?������������������������       �z�G�z�?             @      �?C       D                 �&B@�q�q�?             2@     �?������������������������       �X�<ݚ�?             "@      �?������������������������       ������H�?             "@      �?F       M                    .@�ݏ^���?            �F@     �?G       L                   �*@X�Cc�?             <@     �?H       I                 @33"@�G��l��?             5@      �?������������������������       �      �?              @      �?J       K                 Ь�$@�	j*D�?             *@      �?������������������������       �և���X�?             @      �?������������������������       �r�q��?             @      �?������������������������       �                     @      �?N       O                 ��Y1@������?             1@     �?������������������������       �      �?              @      �?������������������������       ��q�q�?             "@      �?Q       R                    @�nkK�?             7@     �?������������������������       �        
             1@      �?������������������������       �r�q��?             @      �?�t�b��     h�h)h,K ��h.��R�(KKSKK��h\�B0       �|@     @o@     @y@     �V@      @      0@              $@      @      @              @      @      �?      y@     �R@     s@     @Q@     �r@      M@     �n@      D@      0@             �l@      D@      (@             @k@      D@      5@      @      .@      @      @      @     �h@     �@@      :@      @       @              2@      @      (@       @      @      �?     `e@      >@      J@      2@      =@      0@      ;@      "@       @      @      7@       @      $@       @       @               @       @      *@              @      &@      �?      @      @      @     �W@      @      $@       @      @      �?      @      �?     @U@      @      S@      @     �O@       @     �J@              $@       @      @       @      @              *@      �?      "@              M@      d@      @     �[@      @     �X@      @      D@      @      @              B@             �M@      @      (@              $@      @       @      J@     �H@      >@      H@       @      9@       @      *@      �?      "@      �?      @      @      (@      @      @      �?       @      6@      7@      2@      $@      &@      $@      @      �?      @      "@      @      @      �?      @      @              @      *@      �?      @      @      @      6@      �?      1@              @      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�[�.hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKohth)h,K ��h.��R�(KKo��h{�B�         L                    �?@?�p�?�           @�@                                  @>.��Y��?*           `|@      �?                            @�����?             3@        ������������������������       �                      @      �?������������������������       ��eP*L��?             &@      "@       I                    �?u�i-��?           0{@     @                          �;@���e��?           0y@      @                           �?d,���O�?L            �Y@      @	       
                    5@     ��?             0@      @������������������������       ��q�q�?             @     @������������������������       �      �?             $@      �?                        P�@�4���L�?@            �U@      �?������������������������       �և���X�?             @       @                          �:@�P�����?<            �S@                                 �5@L������?8            @R@     .@                           �?&^�)b�?"            �E@     @                        ��Y @��hJ,�?             A@ �������                          �3@������?             1@        ������������������������       ��z�G��?             $@9       ������������������������       �؇���X�?             @8                                 �1@�IєX�?             1@        ������������������������       �      �?             @��������������������������������       �                     *@��������������������������������       ��q�q�?             "@��������������������������������       �                     >@;       ������������������������       �r�q��?             @��������       8                 ��D:@<���n��?�            �r@�������       7                   �L@��r>�?�            `k@             0                    A@��-#���?�            �j@             -                   �*@��cˣ��?_            �b@                                    @����?J            @\@        ������������������������       ���s����?             5@A      !       $                    �?�LQ�1	�?<             W@       "       #                   �<@���@��?            �B@      ������������������������       �\-��p�?             =@�       ������������������������       �      �?              @�       %       &                 �&B@,�+�C�?#            �K@        ������������������������       �                     "@j       '       (                   �<@���}<S�?             G@       ������������������������       �                     =@�       )       ,                   @@@������?             1@       *       +                   �?@�q�q�?             (@        ������������������������       ��q�q�?             @$       ������������������������       ��q�q�?             @       ������������������������       �                     @       .       /                     @�?�|�?            �B@        ������������������������       ��8��8��?             (@]       ������������������������       �                     9@�       1       2                     @0�z��?�?$             O@        ������������������������       �                     6@�       3       4                 �?�@�(\����?             D@       ������������������������       �                     8@�       5       6                 pFt @      �?             0@       ������������������������       �ףp=
�?             $@      ������������������������       �                     @�       ������������������������       �����X�?             @`      9       D                    �?�4F����?7            �T@      :       C                   �J@      �?)             P@      ;       B                    �?��WV��?!             J@      <       ?                   �>@X��ʑ��?            �E@       =       >                    ?@�E��ӭ�?             2@      ������������������������       �X�<ݚ�?             "@G       ������������������������       ������H�?             "@      @       A                 0�K@`�Q��?             9@      ������������������������       ����y4F�?	             3@�      ������������������������       ��q�q�?             @�      ������������������������       ��<ݚ�?             "@8       ������������������������       ��8��8��?             (@8      E       H                     �?�����H�?             2@      F       G                    �?"pc�
�?
             &@       ������������������������       �                     @,      ������������������������       �����X�?             @�      ������������������������       �                     @�       J       K                    �?      �?             @@        ������������������������       �z�G�z�?             @v      ������������������������       �                     ;@�      M       Z                   �2@�+��0��?�             p@       N       Q                     @�ݜ����?"            �M@       O       P                    @�t����?             1@       ������������������������       �����X�?             @�      ������������������������       �                     $@�       R       W                 ��*4@�ՙ/�?             E@      S       V                    �?��
ц��?             :@      T       U                   �0@b�2�tk�?             2@       ������������������������       �և���X�?             @g      ������������������������       ����!pc�?             &@�       ������������������������       �      �?              @y       X       Y                    @      �?             0@        ������������������������       �      �?              @�       ������������������������       �                      @        [       `                     @�y�bm�?y            �h@       \       _                 03[=@�Μ�5�?D            �[@        ]       ^                 `ff:@ �q�q�?             H@       ������������������������       �                     D@        ������������������������       �      �?              @        ������������������������       �        &            �O@        a       b                    �?d�
��?5             V@        ������������������������       ����B���?             :@        c       d                   �@�BE����?%             O@        ������������������������       ������H�?             "@        e       j                    �?�c�����?             �J@        f       i                 `f�%@�eP*L��?             6@       g       h                   @"@z�G�z�?
             .@       ������������������������       �ףp=
�?             $@        ������������������������       ����Q��?             @        ������������������������       �                     @        k       n                 ��1@��a�n`�?             ?@        l       m                   @.@      �?	             (@       ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �        	             3@        �t�bh�h)h,K ��h.��R�(KKoKK��h\�B�       �{@     �p@      w@     �U@      @      *@               @      @      @     �v@     @R@     �t@      R@      S@      :@      @      "@       @      @      @      @     @Q@      1@      @      @     �P@      *@     @P@       @     �A@       @      =@      @      *@      @      @      @      @      �?      0@      �?      @      �?      *@              @      @      >@              �?      @     �o@      G@     �h@      4@     @h@      2@     �`@      1@     @X@      0@      1@      @      T@      (@      =@       @      9@      @      @      @     �I@      @      "@              E@      @      =@              *@      @       @      @      @       @      @       @      @              B@      �?      &@      �?      9@             �N@      �?      6@             �C@      �?      8@              .@      �?      "@      �?      @              @       @      L@      :@      D@      8@      =@      7@      6@      5@      @      *@      @      @      �?       @      1@       @      .@      @       @      @      @       @      &@      �?      0@       @      "@       @      @              @       @      @              ?@      �?      @      �?      ;@              S@     �f@      <@      ?@       @      .@       @      @              $@      :@      0@      (@      ,@      &@      @      @      @       @      @      �?      @      ,@       @      @       @       @              H@     �b@       @     @[@       @      G@              D@       @      @             �O@      G@      E@      @      5@     �D@      5@      �?       @      D@      *@      (@      $@      (@      @      "@      �?      @       @              @      <@      @      "@      @      @              @      @      3@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��=hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKohth)h,K ��h.��R�(KKo��h{�B�         (                     @�)�>_M�?�           @�@                                   �?`՟�G��?�            `s@     �?                           (@�4��`��?q            `f@      @@������������������������       �        	             *@      �?                          �M@4�{Y���?h            �d@     �?                            �?8�Z$���?a            �c@      @       
                   �;@��Sݭg�?0            �S@      4@       	                 Ј@S@�q�q�?             (@      @������������������������       ��q�q�?             @      @������������������������       �      �?             @                                `f�B@F.< ?�?(            �P@      @                           =@�c�Α�?             =@                                ���=@�n_Y�K�?	             *@        ������������������������       �z�G�z�?             @       @������������������������       �      �?              @      5@                        ��:@     ��?             0@       @������������������������       �                     @Z                              ���<@���!pc�?	             &@       ������������������������       ����Q��?             @�      ������������������������       �r�q��?             @w                               x#J@$G$n��?            �B@       ������������������������       �                     (@�                                �D@z�G�z�?             9@       ������������������������       �X�<ݚ�?             "@�                              03�S@      �?             0@       ������������������������       �r�q��?             @c      ������������������������       �                     $@                                �*@�7��?1            �S@      ������������������������       �$�q-�?!             J@�      ������������������������       �                     :@(      ������������������������       ����Q��?             $@V              '                    �?@��A1ʞ?P            ``@      !       &                   �6@����?�?6            �V@       "       #                    �?�X�<ݺ?             B@       ������������������������       �                     $@�       $       %                   �;@$�q-�?             :@        ������������������������       �      �?             @v       ������������������������       �        
             6@j       ������������������������       �        #             K@�       ������������������������       �                    �D@�       )       V                    �?!��)��?�             y@       *       =                 �?�@PN��T'�?�            �p@        +       <                    �?������?X             b@       ,       9                 �{@�#-���?S            �a@       -       2                    �?���z�k�?<            �Y@        .       1                   �=@H%u��?             I@       /       0                   �:@�MI8d�?            �B@        ������������������������       ��<ݚ�?             "@�       ������������������������       �؇���X�?             <@A       ������������������������       �                     *@�       3       8                 �?$@0��_��?!            �J@       4       7                   �:@������?            �D@        5       6                    7@�KM�]�?             3@       ������������������������       �                     ,@      ������������������������       ����Q��?             @�       ������������������������       �                     6@`      ������������������������       �      �?             (@:      :       ;                   �<@�?�|�?            �B@      ������������������������       �                     <@?      ������������������������       ������H�?             "@I      ������������������������       �z�G�z�?             @7      >       ?                 @3�@��n��?Y            @_@        ������������������������       ��q�q�?             (@      @       Q                    �? ��(��?S            @\@      A       B                    �?�ݜ�?;            �S@       ������������������������       ����Q��?             @�      C       P                    �?����1�?7            @R@       D       O                 �T)D@Xny��?.            �N@      E       N                   �>@@4և���?)             L@      F       M                    (@dP-���?!            �G@      G       J                 ��) @�����?             E@       H       I                   �5@�X�<ݺ?             2@       ������������������������       �      �?             @�       ������������������������       �        	             ,@�       K       L                 ���!@      �?             8@       ������������������������       �z�G�z�?             $@�      ������������������������       �@4և���?             ,@�      ������������������������       �                     @�      ������������������������       �                     "@�      ������������������������       ����Q��?             @�      ������������������������       �        	             (@�       R       U                    �?����X�?            �A@      S       T                    0@�n_Y�K�?             :@       ������������������������       ��q�q�?             .@%      ������������������������       �        	             &@g      ������������������������       �                     "@�       W       `                   �7@�'�=z��?F            �`@        X       _                 `f7@���!pc�?            �K@       Y       Z                    @�X���?             F@        ������������������������       ��q�q�?             (@        [       \                    �?     ��?             @@        ������������������������       ��8��8��?             (@        ]       ^                   �5@�z�G��?             4@       ������������������������       ��q�q�?             (@        ������������������������       �      �?              @        ������������������������       �                     &@        a       n                    @���|���?*            @S@       b       m                 03�7@�Y�R_�?&            �Q@       c       f                    �?�<ݚ�?!            �O@        d       e                    �?ףp=
�?             >@       ������������������������       ������H�?
             2@        ������������������������       ��8��8��?             (@        g       j                 P��$@�q�q�?            �@@       h       i                   �=@�q�q�?	             .@       ������������������������       �և���X�?             @        ������������������������       �      �?              @        k       l                    =@�X�<ݺ?             2@        ������������������������       �                     @        ������������������������       ��C��2(�?             &@        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KKoKK��h\�B�       `{@      q@     �a@     @e@     @a@     �D@              *@     @a@      <@     �`@      8@      M@      4@      @      @       @      @      @      @     �J@      *@      5@       @       @      @      @      �?      @      @      *@      @      @               @      @      @       @      @      �?      @@      @      (@              4@      @      @      @      .@      �?      @      �?      $@             �R@      @      H@      @      :@              @      @       @      `@       @      V@       @      A@              $@       @      8@       @       @              6@              K@             �D@     �r@      Z@     �l@      D@     �`@      *@      `@      (@      W@      &@      F@      @      ?@      @      @       @      8@      @      *@              H@      @     �C@       @      1@       @      ,@              @       @      6@              "@      @      B@      �?      <@               @      �?      @      �?     �X@      ;@      @      @     @W@      4@      Q@      $@       @      @     �P@      @      K@      @      J@      @     �E@      @      C@      @      1@      �?      @      �?      ,@              5@      @       @       @      *@      �?      @              "@               @      @      (@              9@      $@      0@      $@      @      $@      &@              "@              Q@      P@      D@      .@      =@      .@      @       @      9@      @      &@      �?      ,@      @       @      @      @       @      &@              <@     �H@      6@     �H@      ,@     �H@      @      ;@       @      0@      �?      &@      &@      6@      $@      @      @      @      @      �?      �?      1@              @      �?      $@       @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��(hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK
hsKmhth)h,K ��h.��R�(KKm��h{�B@         "                 `f�$@(����7�?�           @�@                                   �?�'�`d�?�            �p@     @                          �<@�'����?�             j@     5@                          �;@�1h�'��?b            `b@      .@                           �?H%u��?/            �R@     @       	                 ���@�����?'            �O@      �?                           �?      �?             0@      "@������������������������       ��<ݚ�?             "@        ������������������������       �����X�?             @      @
                           �?`�q�0ܴ?            �G@      �?������������������������       �z�G�z�?             @       @                          �5@�Ń��̧?             E@                                 �@���7�?             6@     �[@������������������������       �؇���X�?             @      B@������������������������       �        	             .@       @������������������������       �                     4@      *@������������������������       �      �?             (@Z                                 �?�X�<ݺ?3             R@       ������������������������       �H%u��?             9@�                              �?$@`Ql�R�?!            �G@                                  @�X�<ݺ?             2@      ������������������������       �                     ,@�      ������������������������       �      �?             @�      ������������������������       �                     =@�                                �=@��a�n`�?*             O@       ������������������������       �      �?              @c                              �&B@r�q��?&             K@       ������������������������       �                     6@      ������������������������       �     ��?             @@�                              ��@\�����?!            �K@       ������������������������       ���s����?             5@V              !                   �>@ҳ�wY;�?             A@      ������������������������       ��	j*D�?             :@3      ������������������������       �      �?              @A      #       6                    �?~h����?            |@        $       1                    �?$�ݏ^��?9            �V@       %       ,                     �?r�q��?             H@       &       +                    �?���>4��?             <@       '       (                 `f�B@�ՙ/�?             5@        ������������������������       ��q�q�?             @�       )       *                 `��W@������?	             .@        ������������������������       �                     @�       ������������������������       ����Q��?             $@$       ������������������������       �                     @       -       0                     @��Q��?             4@       .       /                    �?"pc�
�?             &@        ������������������������       �      �?             @]       ������������������������       �                     @�       ������������������������       �X�<ݚ�?             "@A       2       3                     @@4և���?             E@       ������������������������       �                     <@�       4       5                   �"@d}h���?	             ,@        ������������������������       �                      @�       ������������������������       �      �?             @      7       V                     @�gS��l�?�            `v@       8       O                    �?�ݏ^���?�             l@      9       :                    $@�������?O            �`@       ������������������������       �                     @;      ;       H                     �?�J�4�?J            @_@       <       E                    �?�k�'7��?$            �L@      =       D                   �J@x�����?            �C@      >       A                   @>@`�Q��?             9@        ?       @                    D@d}h���?             ,@       ������������������������       ������H�?             "@!      ������������������������       ����Q��?             @�      B       C                   �@@�eP*L��?	             &@       ������������������������       �z�G�z�?             @8       ������������������������       �r�q��?             @8      ������������������������       �                     ,@      F       G                    �?�����H�?             2@       ������������������������       �                      @,      ������������������������       �z�G�z�?             $@�      I       N                    �?��hJ,�?&             Q@       J       M                   �*@�+$�jP�?              K@       K       L                   �;@�<ݚ�?            �F@       ������������������������       �        
             2@�      ������������������������       ���}*_��?             ;@�      ������������������������       �                     "@�      ������������������������       �                     ,@�      P       U                   �;@ rpa�?=            @W@       Q       T                   �8@؇���X�?            �A@       R       S                   �4@h�����?             <@       ������������������������       �      �?             @-      ������������������������       �                     8@%      ������������������������       �և���X�?             @g      ������������������������       �        $             M@�       W       X                 0S�*@4;����?Q            �`@        ������������������������       �                     (@}       Y       d                    �?�e+��?L            @^@       Z       _                 ��T?@$G$n��?-            �R@       [       \                    )@�C��2(�?            �K@        ������������������������       �����X�?             ,@        ]       ^                    �?��Y��]�?            �D@        ������������������������       �      �?              @        ������������������������       �                    �@@        `       c                    @�d�����?             3@       a       b                 0�H@�eP*L��?	             &@        ������������������������       ��q�q�?             @        ������������������������       ����Q��?             @        ������������������������       �                      @        e       f                    �?֭��F?�?            �G@        ������������������������       �                     @        g       h                    �?��i#[�?             E@        ������������������������       �և���X�?             ,@        i       l                    @      �?             <@       j       k                 �̼6@�S����?             3@        ������������������������       �      �?             @        ������������������������       �        	             *@        ������������������������       �X�<ݚ�?             "@        �t�bh�h)h,K ��h.��R�(KKmKK��h\�B�       �{@      q@      j@      L@     �f@      ;@     �`@      *@     �P@      "@     �L@      @      (@      @      @       @      @       @     �F@       @      @      �?     �D@      �?      5@      �?      @      �?      .@              4@              "@      @      Q@      @      6@      @      G@      �?      1@      �?      ,@              @      �?      =@              H@      ,@      @      @     �F@      "@      6@              7@      "@      :@      =@      @      1@      6@      (@      2@       @      @      @      m@      k@      =@     �N@      :@      6@      *@      .@      *@       @       @      @      &@      @      @              @      @              @      *@      @      "@       @       @       @      @              @      @      @     �C@              <@      @      &@               @      @      @     `i@     `c@     �[@     �\@     @Z@      ;@              @     @Z@      4@     �G@      $@      ?@       @      1@       @      &@      @       @      �?      @       @      @      @      �?      @      @      �?      ,@              0@       @       @               @       @      M@      $@      F@      $@     �A@      $@      2@              1@      $@      "@              ,@              @      V@      @      >@      �?      ;@      �?      @              8@      @      @              M@     @W@      D@              (@     @W@      <@      P@      $@      I@      @      $@      @      D@      �?      @      �?     �@@              ,@      @      @      @      @       @       @      @       @              =@      2@              @      =@      *@       @      @      5@      @      0@      @      @      @      *@              @      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ���~hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKchth)h,K ��h.��R�(KKc��h{�B�                             @�6��l�?�           @�@                                   @�θ�?            �C@      @                           �?�g�y��?             ?@       ������������������������       �                     5@0�G��  ������������������������       �ףp=
�?             $@      �?������������������������       �                      @      @       J                    �?b�h�{��?�           �@     @       G                   �K@j�q����?            |@     `@	                           �?ް� ��?
           �z@      8@
                         A7@�(�Tw��?,            �S@    �D@                        �y�#@X�Cc�?             E@     (@                          �:@d}h���?             <@       @������������������������       ����Q��?             @       @                           ?@�LQ�1	�?             7@       ������������������������       �r�q��?
             2@      �?������������������������       �                     @      4@                          �8@X�Cc�?             ,@       ������������������������       �      �?              @�      ������������������������       ��q�q�?             @�                                 �?tk~X��?             B@                              �D�G@      �?             8@       ������������������������       �                      @�                                �;@      �?	             0@      ������������������������       �      �?              @�      ������������������������       �      �?              @�      ������������������������       ��8��8��?             (@c             8                 ��D:@؇���X�?�            �u@             5                   �*@4z:V��?�            �q@                                �0@�Y��$�?�            �l@       ������������������������       �և���X�?             @(             "                   �7@��(�2Y�?�            �k@               !                    �? �Jj�G�?#            �K@      ������������������������       �                    �G@3      ������������������������       �      �?              @A      #       4                   @F@~n��W��?i            �d@       $       %                     �?z���=��?a            @c@        ������������������������       �                     @v       &       1                 `fF)@��H�&p�?\            �b@       '       ,                 @3�@D|U��@�?T            �`@       (       +                    �?�[$�G�?;            �X@        )       *                  s�@�LQ�1	�?             7@        ������������������������       �                     @�       ������������������������       �@�0�!��?
             1@$       ������������������������       �DE��2{�?-            �R@       -       .                     @������?             B@        ������������������������       �                     @-       /       0                 @Q!@�g�y��?             ?@       ������������������������       �                     8@�       ������������������������       �؇���X�?             @A       2       3                   �;@���Q��?             .@        ������������������������       �                      @�       ������������������������       �؇���X�?             @�       ������������������������       �                     *@�       6       7                    �?�h����?!             L@       ������������������������       �r�q��?             @�       ������������������������       �                     I@`      9       B                     �?R=6�z�?-            @P@      :       ?                    �?�J��%�?            �H@      ;       <                   �@@h+�v:�?             A@      ������������������������       �      �?             0@I      =       >                 `f�<@      �?
             2@       ������������������������       �      �?              @G       ������������������������       �z�G�z�?             $@      @       A                   �C@z�G�z�?
             .@       ������������������������       �      �?              @�      ������������������������       �                     @�      C       F                    �?     ��?             0@       D       E                    ;@      �?              @       ������������������������       �      �?             @      ������������������������       �      �?             @-      ������������������������       �                      @,      H       I                   �O@8�A�0��?             6@      ������������������������       �     ��?             0@�       ������������������������       �                     @�       K       `                 ���H@� ��Z�?�            �k@      L       ]                 03�;@��Q��?h             d@      M       R                     @�����?Z             a@       N       Q                   �6@�X�<ݺ?$             K@      O       P                   �;@ףp=
�?             >@       ������������������������       ����!pc�?             &@�      ������������������������       �                     3@�       ������������������������       �                     8@      S       X                    �?F~��7�?6            �T@       T       W                    �?؇���X�?             <@      U       V                 ���@؇���X�?             5@       ������������������������       �                     "@�       ������������������������       �      �?             (@y       ������������������������       �؇���X�?             @}       Y       Z                    �?ؓ��M{�?$            �K@       ������������������������       ���S���?             >@        [       \                 ���4@`�Q��?             9@       ������������������������       ���.k���?             1@        ������������������������       �                      @        ^       _                     @��<b���?             7@        ������������������������       �      �?              @        ������������������������       �        	             .@        a       b                    �? ������?&            �O@       ������������������������       �                     �K@        ������������������������       �      �?              @        �t�bh�h)h,K ��h.��R�(KKcKK��h\�B0       0{@     Pq@      "@      >@      �?      >@              5@      �?      "@       @             �z@     �n@     w@     @T@     @v@      R@      L@      6@      ;@      .@      6@      @       @      @      4@      @      .@      @      @              @      "@      @      @       @      @      =@      @      2@      @       @              $@      @      @      @      @      �?      &@      �?     �r@      I@     �o@      ?@     �h@      >@      @      @     `h@      ;@      K@      �?     �G@              @      �?     �a@      :@      `@      :@      @             �^@      :@     �\@      4@     �S@      3@      4@      @      @              ,@      @     �M@      0@     �A@      �?      @              >@      �?      8@              @      �?      "@      @       @              �?      @      *@             �K@      �?      @      �?      I@              G@      3@     �@@      0@      5@      *@      (@      @      "@      "@      �?      @       @       @      (@      @      @      @      @              *@      @      @      @       @       @      @      �?       @              *@      "@      @      "@      @             �L@     �d@      L@      Z@      C@     �X@      @     �I@      @      ;@      @       @              3@              8@     �A@      H@      @      8@      @      2@              "@      @      "@      �?      @      ?@      8@      ,@      0@      1@       @      "@       @       @              2@      @      @      @      .@              �?      O@             �K@      �?      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJCLUhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKghth)h,K ��h.��R�(KKg��h{�B�         .                     @Dl���v�?�           @�@               %                  ��T@d ���T�?�            �s@    @T@                           �?t����?�            �p@     @       	                 ��\+@ޭ�W[��?i            @d@                                  �@@�q��/��?!            �H@     �?������������������������       �                    �@@                                  �B@      �?             0@        ������������������������       �      �?             @      (@������������������������       ��z�G��?             $@     �N@
                           �?4;W!���?H            @\@     @                           @@�7�A�?4             V@      @                           �?�q�q�?             B@        ������������������������       ��eP*L��?             &@      &@                           �? �o_��?             9@    �\@                          �>@      �?	             (@     $@������������������������       ����Q��?             @      �?������������������������       �                     @Z      ������������������������       ��	j*D�?             *@�                              ��$:@D>�Q�?             J@       ������������������������       �        	             .@w                                �G@���"͏�?            �B@                                 �E@�����H�?	             2@       ������������������������       ��<ݚ�?             "@�      ������������������������       �                     "@�      ������������������������       �p�ݯ��?             3@�                                 +@� �	��?             9@       ������������������������       �                     "@                              ���G@      �?             0@      ������������������������       �                     $@�      ������������������������       ��q�q�?             @(             "                    �?�]��?:            �Y@               !                    �?�����?             5@       ������������������������       �����X�?             @3      ������������������������       �                     ,@A      #       $                    6@��Y��]�?.            �T@        ������������������������       ��FVQ&�?            �@@�       ������������������������       �                    �H@v       &       )                    �?f1r��g�?"            �J@       '       (                    �?@4և���?             <@        ������������������������       ����Q��?             @�       ������������������������       �                     7@�       *       -                   @C@�+e�X�?             9@       +       ,                 03�a@R���Q�?             4@       ������������������������       �                     (@       ������������������������       �      �?              @       ������������������������       ����Q��?             @-       /       T                    �?��머��?�            �x@       0       S                 �T�I@��W��?�            �q@       1       L                    �?,T\��?�            �p@       2       G                 ��i @ܷ��?��?�             m@       3       @                   �<@      �?i             f@       4       5                    �?85�}C�?G            �^@        ������������������������       ��S����?             3@�       6       7                   �4@b �57�?;            �Y@       ������������������������       �                     <@�       8       =                   �9@���Lͩ�?.            �R@       9       <                 ��L@�㙢�c�?             7@      :       ;                    7@���|���?	             &@       ������������������������       �      �?             @?      ������������������������       �և���X�?             @I      ������������������������       �                     (@7      >       ?                    �?0G���ջ?             J@        ������������������������       �P���Q�?             4@      ������������������������       �      �?             @@!      A       D                   @@@�<ݚ�?"             K@       B       C                   �?@D�n�3�?             3@      ������������������������       �X�<ݚ�?             "@8       ������������������������       ��z�G��?             $@8      E       F                 �?�@��?^�k�?            �A@      ������������������������       �                     7@-      ������������������������       ��8��8��?             (@,      H       I                 ���"@h�����?"             L@       ������������������������       �                     <@�       J       K                 �&�)@@4և���?             <@        ������������������������       �����X�?             @v      ������������������������       �                     5@�      M       P                    @      �?             B@      N       O                    /@�LQ�1	�?             7@       ������������������������       �      �?              @�      ������������������������       ���S�ۿ?	             .@�      Q       R                    �?$�q-�?	             *@       ������������������������       �                     "@      ������������������������       �      �?             @-      ������������������������       ��q�q�?             (@%      U       d                    @6C�z��?G            �\@      V       c                 ��Y7@�q�Q�?<             X@       W       X                    "@b�2�tk�?8            �V@        ������������������������       �                     @}       Y       Z                    �?j���� �?4            @U@        ������������������������       ��z�G��?             $@        [       b                   �@@L�qA��?/            �R@       \       _                    �?<��¤�?+             Q@        ]       ^                    9@      �?             <@        ������������������������       ��q�q�?             @        ������������������������       ��GN�z�?             6@        `       a                    �?      �?             D@       ������������������������       ��P�*�?             ?@        ������������������������       ��<ݚ�?             "@        ������������������������       �؇���X�?             @        ������������������������       �                     @        e       f                   �6@r�q��?             2@       ������������������������       �      �?              @        ������������������������       �                     $@        �t�bh�h)h,K ��h.��R�(KKgKK��h\�Bp        {@     `q@      a@     �f@      `@      a@      _@      C@     �E@      @     �@@              $@      @      @      @      @      @     @T@      @@     �P@      5@      8@      (@      @      @      2@      @      "@      @       @      @      @              "@      @     �E@      "@      .@              <@      "@      0@       @      @       @      "@              (@      @      ,@      &@              "@      ,@       @      $@              @       @      @     �X@       @      3@       @      @              ,@       @      T@       @      ?@             �H@       @     �F@       @      :@       @      @              7@      @      3@      @      1@              (@      @      @      @       @     �r@      X@     @n@      C@     `m@     �@@      j@      8@     @c@      6@      \@      $@      0@      @      X@      @      <@              Q@      @      3@      @      @      @      @      �?      @      @      (@             �H@      @      3@      �?      >@       @      E@      (@       @      &@      @      @      @      @      A@      �?      7@              &@      �?      K@       @      <@              :@       @      @       @      5@              ;@      "@      .@       @      �?      @      ,@      �?      (@      �?      "@              @      �?      @      @      L@      M@     �D@     �K@     �A@     �K@              @     �A@      I@      @      @      <@     �G@      ;@     �D@      @      5@       @      @      @      1@      4@      4@      *@      2@      @       @      �?      @      @              .@      @      @      @      $@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ���hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKqhth)h,K ��h.��R�(KKq��h{�B@         0                     @#�[5]�?�           @�@               !                    �?�B܎���?�            ps@     ;@                           (@yp3�?s             g@      *@������������������������       �                     @     @                         I>@$�����?n            `f@     @                           �?�=|+g��?D            @\@     @       
                   �@@ףp=
�?7            �V@      ?@       	                    5@���7�?             F@      �?������������������������       �      �?              @      :@������������������������       �������?             B@      3@                            �?*
;&���?             G@      0@������������������������       �      �?	             0@                                   F@r�q��?             >@      @������������������������       ��	j*D�?	             *@                                  �*@�IєX�?
             1@     @������������������������       �ףp=
�?             $@      @������������������������       �                     @Z                                 :@�nkK�?             7@      ������������������������       �@4և���?             ,@�      ������������������������       �                     "@w                                �?@���!pc�?*            �P@       ������������������������       ��<ݚ�?             "@�                                �8@F�t�K��?&            �L@       ������������������������       �                     "@�                                 �?�q�q��?             H@       ������������������������       ��q�q�?	             (@c                                  �?tk~X��?             B@                                 �?�+$�jP�?             ;@       ������������������������       �8�Z$���?             *@�                              ���O@d}h���?	             ,@       ������������������������       ����Q��?             @V      ������������������������       ������H�?             "@J      ������������������������       ��<ݚ�?             "@3      "       %                    6@$Q�q�?O            �_@       #       $                   �;@�r����?             >@        ������������������������       �X�<ݚ�?             "@�       ������������������������       �                     5@v       &       '                    @ �q�q�?=             X@        ������������������������       �z�G�z�?             @�       (       -                    �?x��B�R�?8            �V@       )       ,                    �? �й���?-            @R@        *       +                   �H@�}�+r��?             3@       ������������������������       �                     .@$       ������������������������       �      �?             @       ������������������������       �                     K@       .       /                   �8@�����H�?             2@       ������������������������       �                      @]       ������������������������       �z�G�z�?             $@�       1       6                    @X-�?2�?�            y@        2       5                    �?�g�y��?             ?@       3       4                    �?      �?
             0@        ������������������������       �r�q��?             @�       ������������������������       ��z�G��?             $@�       ������������������������       �������?             .@      7       n                 ��Y7@yp3�?�             w@       8       c                    �?Z]k�Β�?�            �t@      9       V                    �?|���~�?�             q@      :       Q                   @@@$Nz�{�?�             k@      ;       L                   �<@�S-�?j            �d@      <       ?                    �?���;QU�?[            @b@       =       >                    ;@�����H�?             ;@       ������������������������       �      �?             @G       ������������������������       �        	             5@      @       A                 ��Y@�IєX�?N            �]@       ������������������������       �z�G�z�?             $@�      B       G                 @3�@ '��h�?I            @[@      C       F                 ��@0�)AU��?(            �L@        D       E                   �:@���N8�?             5@       ������������������������       �                      @      ������������������������       �$�q-�?	             *@-      ������������������������       �                     B@,      H       K                 ��i @$�q-�?!             J@      I       J                   �3@\-��p�?             =@        ������������������������       �և���X�?             @�       ������������������������       ����7�?             6@v      ������������������������       �                     7@�      M       N                 �?�@����X�?             5@       ������������������������       �r�q��?             @�      O       P                   �>@�q�q�?
             .@       ������������������������       �r�q��?             @�      ������������������������       �X�<ݚ�?             "@�       R       S                 �?�@p���?!             I@      ������������������������       �                     >@-      T       U                 pFt @P���Q�?             4@       ������������������������       �ףp=
�?             $@g      ������������������������       �                     $@�       W       `                    �?F�����?%            �L@       X       [                    �?X��ʑ��?            �E@        Y       Z                 �&B@b�2�tk�?             2@       ������������������������       ��q�q�?             (@        ������������������������       �      �?             @        \       _                 `�X!@� �	��?             9@       ]       ^                  sW@      �?             0@        ������������������������       �      �?              @        ������������������������       �      �?              @        ������������������������       �X�<ݚ�?             "@        a       b                   �;@X�Cc�?             ,@        ������������������������       �؇���X�?             @        ������������������������       �և���X�?             @        d       e                 pf� @�q�q�?#             K@        ������������������������       �      �?             $@        f       g                    ;@v�X��?             F@        ������������������������       ��C��2(�?             &@        h       m                    �?���|���?            �@@       i       l                   @A@���Q��?             9@       j       k                    �?�q�q�?             2@        ������������������������       �                      @        ������������������������       ����Q��?             $@        ������������������������       �և���X�?             @        ������������������������       �      �?              @        o       p                 0�H@���N8�?             E@       ������������������������       �                     @@        ������������������������       �z�G�z�?             $@        �t�bh�h)h,K ��h.��R�(KKqKK��h\�B       �}@     �m@     �c@      c@     �b@      A@              @     �b@      <@     �Y@      $@     @T@      "@      E@       @      @      �?     �A@      �?     �C@      @      ,@       @      9@      @      "@      @      0@      �?      "@      �?      @              6@      �?      *@      �?      "@              H@      2@       @      @      G@      &@      "@             �B@      &@       @      @      =@      @      6@      @      &@       @      &@      @      @       @       @      �?      @       @       @     �]@      @      :@      @      @              5@      @      W@      �?      @      @      V@      �?      R@      �?      2@              .@      �?      @              K@       @      0@               @       @       @     �s@      U@      .@      0@      @      (@      �?      @      @      @      &@      @     �r@      Q@     `p@     �P@     @l@      H@      i@      1@     �b@      0@      a@      $@      8@      @      @      @      5@              \@      @       @       @      Z@      @      L@      �?      4@      �?       @              (@      �?      B@              H@      @      9@      @      @      @      5@      �?      7@              .@      @      @      �?      $@      @      @      �?      @      @     �H@      �?      >@              3@      �?      "@      �?      $@              :@      ?@      5@      6@      @      &@      @       @      @      @      ,@      &@      $@      @      @      @      @       @      @      @      @      "@      �?      @      @      @      B@      2@      @      @      ?@      *@      $@      �?      5@      (@      .@      $@      (@      @       @              @      @      @      @      @       @      D@       @      @@               @       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ"�a,hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKmhth)h,K ��h.��R�(KKm��h{�B@         
                    @�6��l�?�           @�@                                   @�^�����?            �E@�X��                          �%D@��a�n`�?             ?@                                  �?`2U0*��?             9@ ��4    ������������������������       ��C��2(�?             &@        ������������������������       �        	             ,@        ������������������������       ��q�q�?             @               	                    @r�q��?             (@        ������������������������       �                     @      ?@������������������������       ����Q��?             @      @       `                  x#J@`S�as��?�           �@     (@       /                     @Ҷx�Т�?g           @�@      C@                          �;@=���?x             g@      $@                           �?p�v>��?            �G@      @                          �3@     ��?             0@     @������������������������       �                     $@       @������������������������       �      �?             @Z                                 �?�g�y��?             ?@                              �J,@P���Q�?             4@       ������������������������       �r�q��?             @w      ������������������������       �                     ,@n      ������������������������       �                     &@�             $                 `f�:@�#��ؒ�?[            @a@             !                   �I@$)}�~z�?>            �W@                                  �?L������?2            �S@                              `ff:@r�q��?             H@                              ��\+@�7��?            �C@      ������������������������       �                     7@                                �@@      �?
             0@      ������������������������       �z�G�z�?             $@(      ������������������������       �                     @V      ������������������������       ��q�q�?             "@J      ������������������������       �                     ?@3      "       #                   �8@�r����?             .@       ������������������������       ��q�q�?             @�       ������������������������       �                     "@�       %       ,                   �E@�������?             F@       &       +                   �>@�C��2(�?            �@@       '       *                    �?R���Q�?             4@       (       )                   �<@      �?             (@        ������������������������       �����X�?             @�       ������������������������       �z�G�z�?             @�       ������������������������       �                      @$       ������������������������       �                     *@       -       .                   �I@�eP*L��?	             &@        ������������������������       �      �?             @-       ������������������������       ����Q��?             @]       0       _                 ��Y7@�Z{����?�            �v@       1       ^                 `v�5@�ɫ5k��?�            �t@       2       K                    �?R���Q�?�             t@       3       4                   �0@��L9���?�            `n@        ������������������������       ��q�q�?             (@�       5       H                 @3�@�s�c���?�            �l@       6       G                 �?�@x�5?,R�?Z             b@      7       :                    �?A5Xo�?R            ``@        8       9                   @@�n`���?             ?@      ������������������������       ��+$�jP�?             ;@:      ������������������������       �      �?             @;      ;       F                    �?HP�s��?@             Y@      <       C                   �?@���.�6�?<             W@      =       >                 ��@�nkK�?/            @Q@       ������������������������       �z�G�z�?             @G       ?       B                   �;@      �?+             P@      @       A                   �9@�IєX�?             A@      ������������������������       �h�����?             <@�      ������������������������       �r�q��?             @�      ������������������������       �                     >@8       D       E                   �@@�LQ�1	�?             7@       ������������������������       ����!pc�?             &@      ������������������������       �                     (@-      ������������������������       �      �?              @,      ������������������������       ��n_Y�K�?             *@�      I       J                    �?X��%�?:            �U@        ������������������������       �      �?             @�       ������������������������       ���`qM|�?6            �T@v      L       U                 @3�@��j��?9            @S@       M       R                    �?      �?             D@      N       O                    9@      �?             4@       ������������������������       �      �?             @�      P       Q                 ���@      �?             0@       ������������������������       �      �?             @�       ������������������������       �      �?             (@      S       T                   �5@      �?             4@       ������������������������       ��z�G��?             $@%      ������������������������       �z�G�z�?             $@g      V       [                    .@^H���+�?            �B@       W       Z                   �=@�㙢�c�?             7@       X       Y                    �?�KM�]�?             3@       ������������������������       ���S�ۿ?             .@�       ������������������������       �      �?             @        ������������������������       �      �?             @        \       ]                 03�1@X�Cc�?             ,@       ������������������������       �                      @        ������������������������       �r�q��?             @        ������������������������       ������H�?             "@        ������������������������       �                     C@        a       h                    �?�(�Tw��?L            @]@        b       g                 `��`@��c:�?             G@       c       f                   �H@      �?             A@       d       e                    @@���Q��?             9@       ������������������������       ����!pc�?	             &@        ������������������������       �؇���X�?             ,@        ������������������������       ��<ݚ�?             "@        ������������������������       �r�q��?             (@        i       j                    �?@�j;��?/            �Q@       ������������������������       �        #            �K@        k       l                    @      �?             0@       ������������������������       �"pc�
�?             &@        ������������������������       �z�G�z�?             @        �t�bh�h)h,K ��h.��R�(KKmKK��h\�B�       0{@     Pq@      *@      >@      @      <@      �?      8@      �?      $@              ,@       @      @      $@       @      @              @       @     `z@     �n@     Px@     `d@     �Y@     �T@      ,@     �@@      *@      @      $@              @      @      �?      >@      �?      3@      �?      @              ,@              &@      V@      I@     �J@     �D@      D@     �C@      D@       @     �B@       @      7@              ,@       @       @       @      @              @      @              ?@      *@       @      @       @      "@             �A@      "@      >@      @      1@      @      "@      @      @       @      @      �?       @              *@              @      @      @      @       @      @     �q@      T@      o@      T@      o@      R@     �j@      =@      @      @     �i@      8@     @_@      3@     @]@      ,@      9@      @      6@      @      @      �?      W@       @     �U@      @     �P@      @      @      �?      O@       @      @@       @      ;@      �?      @      �?      >@              4@      @       @      @      (@              @       @       @      @     �T@      @      @      �?     �S@      @      A@     �E@      $@      >@      @      .@      �?      @      @      (@      �?      @      @      "@      @      .@      @      @       @       @      8@      *@      3@      @      1@       @      ,@      �?      @      �?       @       @      @      "@               @      @      �?      �?       @      C@             �@@      U@      ;@      3@      1@      1@      $@      .@       @      @       @      (@      @       @      $@       @      @     @P@             �K@      @      $@       @      "@      @      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�8�hhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKohth)h,K ��h.��R�(KKo��h{�B�         Z                  x#J@���x�W�?�           @�@                               `f#@�������?x           p�@      �?                          �0@f?�ϼ��?�            `p@        ������������������������       �z�G�z�?             $@      �?                           �?0,Tg��?�            �o@     @                           �?�:�H:�?�            @k@    �D@                           �?�������?�            `i@                                  @@      �?             <@     @	       
                 ���@����X�?
             5@      @������������������������       �z�G�z�?             .@      V@������������������������       �      �?             @      @������������������������       �؇���X�?             @       @                            @p}"����?r            �e@      @������������������������       �                     *@     �P@                        ���@|E+�	��?k            @d@      $@������������������������       �        
             *@      @                        ��}@�
�@c�?a            �b@       ������������������������       ��<ݚ�?             "@�      ������������������������       ����2���?Z            �a@�      ������������������������       ��r����?             .@w                                �5@      �?             A@       ������������������������       �      �?              @�                                 �?�n_Y�K�?             :@       ������������������������       �ףp=
�?             $@�                                �;@     ��?             0@       ������������������������       �      �?              @c      ������������������������       �      �?              @             I                    �?�2�?�            �t@             H                 �D C@Pu�����?�             h@             %                    �?(��a��?t            �e@                                  �8@X�<ݚ�?             ;@       ������������������������       �      �?              @J      !       $                   �=@�����?             3@      "       #                 м;4@"pc�
�?	             &@      ������������������������       �����X�?             @�       ������������������������       �                     @�       ������������������������       �      �?              @v       &       /                     �?� ��fd�?c            @b@        '       .                    K@��}*_��?             ;@       (       -                   �>@�\��N��?             3@       )       *                 03k:@��
ц��?             *@        ������������������������       ����Q��?             @�       +       ,                 `f�;@      �?              @        ������������������������       �      �?             @       ������������������������       �      �?             @       ������������������������       ��q�q�?             @-       ������������������������       �      �?              @]       0       A                    �?p�5�9��?M            �]@       1       2                    �?H��?"�?2             U@        ������������������������       �      �?             @�       3       :                    ?@��-�=��?.            �S@        4       9                    �?������?             B@       5       8                     @h�����?             <@       6       7                    5@���N8�?             5@       ������������������������       �؇���X�?             @�       ������������������������       �                     ,@`      ������������������������       �                     @:      ������������������������       �                      @;      ;       >                   �*@r�q��?             E@       <       =                 `f�)@���N8�?             5@      ������������������������       �"pc�
�?             &@7      ������������������������       ��z�G��?             $@G       ?       @                    C@�����?             5@       ������������������������       �      �?              @!      ������������������������       �                     *@�      B       C                 @3�4@^������?            �A@       ������������������������       �����X�?             ,@8       D       G                    �?�����?             5@      E       F                   �;@�8��8��?
             (@       ������������������������       �z�G�z�?             @-      ������������������������       �                     @,      ������������������������       ������H�?             "@�      ������������������������       �                     4@�       J       K                     @f.i��n�?S            �`@        ������������������������       �        &             P@v      L       O                    �?DX�\��?-            �Q@       M       N                 �?�-@ҳ�wY;�?             1@       ������������������������       �                     @�      ������������������������       �                     &@�      P       Q                    @�q�q�?!             K@       ������������������������       ��q�q�?             (@�       R       S                    -@0,Tg��?             E@       ������������������������       �                     @-      T       Y                 ���4@">�֕�?            �A@      U       V                    �?
;&����?             7@       ������������������������       �      �?             $@�       W       X                 @3�/@��
ц��?	             *@       ������������������������       �      �?              @}       ������������������������       ����Q��?             @�       ������������������������       �                     (@        [       j                 03?U@��6}��?H            �^@       \       _                   �;@�7�֥��?'            @P@        ]       ^                 ���Q@�IєX�?             1@       ������������������������       �                     (@        ������������������������       �z�G�z�?             @        `       c                    �?�q���?             H@        a       b                    �?����X�?             ,@        ������������������������       �X�<ݚ�?             "@        ������������������������       �                     @        d       g                    �?�ʻ����?             A@       e       f                   �D@���y4F�?             3@       ������������������������       �X�<ݚ�?             "@        ������������������������       �                     $@        h       i                   �A@������?	             .@        ������������������������       ��q�q�?             @        ������������������������       �                     "@        k       n                    �?Ԫ2��?!            �L@       l       m                    �?8��8���?             H@        ������������������������       ��eP*L��?             &@        ������������������������       �                    �B@        ������������������������       ��q�q�?             "@        �t�b��     h�h)h,K ��h.��R�(KKoKK��h\�B�       P{@     0q@     Py@      g@     �j@     �G@       @       @     �j@     �C@     �h@      6@     �f@      4@      5@      @      .@      @      (@      @      @      @      @      �?     @d@      *@      *@             �b@      *@      *@              a@      *@      @       @      `@      &@      *@       @      1@      1@      @      �?      $@      0@      �?      "@      "@      @       @      @      @      �?     �g@     @a@     �b@     �F@      `@     �F@      .@      (@       @      @      *@      @      "@       @      @       @      @              @      @     @\@     �@@      1@      $@      $@      "@      @      @       @      @      @      @       @       @       @       @      @       @      @      �?      X@      7@     @R@      &@      @      @     �Q@       @     �A@      �?      ;@      �?      4@      �?      @      �?      ,@              @               @             �A@      @      0@      @      "@       @      @      @      3@       @      @       @      *@              7@      (@      @      $@      3@       @      &@      �?      @      �?      @               @      �?      4@              E@     @W@              P@      E@      =@      @      &@      @                      &@      B@      2@      @      @      ?@      &@      @              8@      &@      (@      &@      @      @      @      @      @      @      @       @      (@              @@     �V@      8@     �D@      �?      0@              (@      �?      @      7@      9@      @      $@      @      @              @      3@      .@      .@      @      @      @      $@              @      &@      @       @              "@       @     �H@      @     �E@      @      @             �B@      @      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJP�dhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK	hsKWhth)h,K ��h.��R�(KKW��h{�B�         @                    �?~�Я��?�           @�@              '                 03�9@ꀕ<u�?%           �}@     @@       &                    �?0���)��?�            �t@      @                        ��y @d��C��?�            `s@     @                        �?�@�t�~U�?o            �f@      @                          �9@@4և���?Q            �_@      "@                          �3@���@��?            �B@     @a@������������������������       �                     @      @	                        �Y�@      �?             @@        
                        ���@     ��?	             0@      @������������������������       �؇���X�?             @        ������������������������       ��q�q�?             "@      T@                          �5@      �?             0@      @������������������������       �z�G�z�?             @      @������������������������       �                     &@      @                        ��@ }�Я��?8            @V@      @������������������������       �        )             P@Z                                 �?`2U0*��?             9@       ������������������������       �z�G�z�?             @�      ������������������������       �                     4@w                              @3�@x��}�?            �K@                                 �?@�eP*L��?             &@       ������������������������       �և���X�?             @�      ������������������������       �      �?             @�      ������������������������       �fP*L��?             F@�                                 �?H*C�|F�?L             `@                                  �?�S����?             3@      ������������������������       �r�q��?             (@      ������������������������       �؇���X�?             @�             !                     @h㱪��?@            �[@                                  �;@�X�<ݺ?              K@       ������������������������       �                     :@J      ������������������������       � �Cc}�?             <@3      "       %                 ���#@�h����?              L@      #       $                   �<@XB���?             =@       ������������������������       �                     .@�       ������������������������       �@4և���?             ,@v       ������������������������       �                     ;@j       ������������������������       ��eP*L��?             6@�       (       ?                    @ޚ)�?Z             b@       )       0                   �>@�����?L            �_@        *       /                   �J@      �?             M@       +       .                    �?nM`����?             G@       ,       -                    ?@����X�?            �A@        ������������������������       �z�G�z�?             $@       ������������������������       �HP�s��?             9@-       ������������������������       ����|���?             &@]       ������������������������       �                     (@�       1       2                   �A@8����?-            @Q@        ������������������������       �                     &@�       3       4                   �9@o����?'             M@        ������������������������       ��C��2(�?             &@�       5       <                    D@�[�IJ�?            �G@       6       9                 `f�N@|��?���?             ;@       7       8                    �?z�G�z�?             $@        ������������������������       �r�q��?             @`      ������������������������       �      �?             @:      :       ;                   �@@ҳ�wY;�?
             1@      ������������������������       �ףp=
�?             $@?      ������������������������       �����X�?             @I      =       >                   �G@�z�G��?             4@       ������������������������       �                     @G       ������������������������       �և���X�?             ,@      ������������������������       �                     1@!      A       H                     @��mo*�?�            �m@      B       C                     �?��G^�C�?S            @`@      ������������������������       �        0            �S@8       D       G                   �8@���J��?#            �I@       E       F                   �+@�}�+r��?             3@       ������������������������       �؇���X�?             @-      ������������������������       �                     (@,      ������������������������       �                     @@�      I       R                    �?��U��?B            �Z@       J       O                   �9@����"�?&             M@        K       L                    �?      �?             @@       ������������������������       �      �?             @�      M       N                    �?���>4��?             <@       ������������������������       �      �?             @�      ������������������������       ��eP*L��?             6@�      P       Q                    �?�θ�?             :@      ������������������������       ������H�?             2@�       ������������������������       �      �?              @      S       V                    �?     ��?             H@      T       U                    .@     ��?             @@       ������������������������       �ףp=
�?             $@g      ������������������������       ����|���?             6@�       ������������������������       �        
             0@y       �t�bh�h)h,K ��h.��R�(KKWKK��h\�Bp       �{@     �p@     0x@     @V@     Pr@     �C@     �q@      =@     �c@      6@     @]@      "@      =@       @      @              8@       @      "@      @      @      �?      @      @      .@      �?      @      �?      &@              V@      �?      P@              8@      �?      @      �?      4@              E@      *@      @      @      @      @       @       @     �B@      @     �^@      @      0@      @      $@       @      @      �?     �Z@      @     �I@      @      :@              9@      @     �K@      �?      <@      �?      .@              *@      �?      ;@              (@      $@     �W@      I@     @S@      I@      =@      =@      1@      =@      $@      9@       @       @       @      7@      @      @      (@              H@      5@      &@             �B@      5@      $@      �?      ;@      4@      *@      ,@       @       @      �?      @      �?      @      &@      @      "@      �?       @      @      ,@      @      @               @      @      1@              L@     �f@      �?      `@             �S@      �?      I@      �?      2@      �?      @              (@              @@     �K@     �I@      6@      B@      0@      0@      �?      @      .@      *@      @      @      (@      $@      @      4@       @      0@      @      @     �@@      .@      1@      .@      "@      �?       @      ,@      0@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�g?BhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKkhth)h,K ��h.��R�(KKk��h{�B�         J                    �?@?�p�?�           @�@              E                    �?@h���?$           `|@                                  @(Z�oh�?           �z@      �?������������������������       �                      @               D                   �M@��a,3�?
           0z@              1                 `ff:@"����U�?           @y@      @       0                   �C@�? Da�?�            �s@      @                        ��y @t�6Z���?�            0q@       	                          �>@���Y�*�?k            �f@       
                           �?13 O��?]            �c@     "@                          �;@��)�c{�?X             c@       @������������������������       �>���Rp�?"             M@      7@                          �<@heu+��?6            �W@     �?                           �?(�s���?0             U@                                 s�@      �?             @@      @                        ���@��S�ۿ?
             .@       @������������������������       �                     @��%�����������������������������       ��C��2(�?             &@.������������������������������       �@�0�!��?             1@w��h�7�                        �?�@ pƵHP�?             J@>\��9s������������������������       �                     B@,������������������������������       �      �?	             0@�iK�Xk"g������������������������       �z�G�z�?             $@�)nɨp������������������������       ��q�q�?             @���y��_                           �?�LQ�1	�?             7@ ��q K������������������������       �                     @2��",}V�������������������������       ���.k���?
             1@+���(��       !                   �9@��8��)�??            �W@ J�EV���                           �3@��Y��]�?            �D@ Z���                           &@      �?
             0@�9(?E�������������������������       �      �?              @��A��������������������������       �                      @rI�L��Pv������������������������       �                     9@3      "       /                    �?f1r��g�?(            �J@      #       &                 `fF)@"pc�
�?#             F@        $       %                   �=@      �?             0@        ������������������������       �      �?              @v       ������������������������       �                      @j       '       *                 �R,@d}h���?             <@        (       )                    @@      �?              @        ������������������������       �      �?             @�       ������������������������       �      �?             @�       +       ,                    �?R���Q�?             4@        ������������������������       �      �?             @       -       .                 039@      �?             0@       ������������������������       �                      @-       ������������������������       �      �?              @]       ������������������������       �                     "@�       ������������������������       �                     D@A       2       ?                    �?:��?=            @V@       3       >                    �?և���X�?(             L@       4       =                      @X��ʑ��?            �E@       5       <                   �G@��%��?            �B@       6       9                    �?��>4և�?             <@       7       8                 `f�C@      �?             $@        ������������������������       ����Q��?             @`      ������������������������       ����Q��?             @:      :       ;                   �>@�q�q�?             2@       ������������������������       �      �?              @?      ������������������������       �ףp=
�?             $@I      ������������������������       ��q�q�?             "@7      ������������������������       �r�q��?             @G       ������������������������       �8�Z$���?
             *@      @       C                   @C@"pc�
�?            �@@      A       B                 `fFJ@���!pc�?             6@       ������������������������       �                     @�      ������������������������       ����Q��?	             .@8       ������������������������       �                     &@8      ������������������������       ���S���?	             .@      F       G                 ��T?@�>����?             ;@      ������������������������       �                     2@,      H       I                     @�<ݚ�?             "@       ������������������������       �      �?             @�       ������������������������       �                     @�       K       T                     @�l]G���?�             p@      L       S                   �;@     p�?W             `@       M       N                    �?Du9iH��?            �E@       ������������������������       �                     .@�      O       P                    �? �Cc}�?             <@       ������������������������       ��<ݚ�?             "@�      Q       R                   0G@�}�+r��?             3@       ������������������������       �                     *@      ������������������������       �r�q��?             @-      ������������������������       �        8            @U@%      U       Z                 pF @^��>�b�?R            @`@       V       W                   �3@���"͏�?            �B@        ������������������������       �X�<ݚ�?             "@y       X       Y                    8@�>4և��?             <@        ������������������������       �                     @�       ������������������������       ���<b���?             7@        [       f                 ���4@���U��?9            @W@       \       c                    �?>n�T��?'             M@       ]       b                    .@�q�q�?             E@       ^       a                  �#@ȵHPS!�?             :@       _       `                   #@P���Q�?             4@       ������������������������       �                     &@        ������������������������       ������H�?             "@        ������������������������       ��q�q�?             @        ������������������������       �     ��?	             0@        d       e                 �&2.@     ��?             0@       ������������������������       ��q�q�?	             (@        ������������������������       �                     @        g       j                    @؇���X�?            �A@       h       i                    �?�nkK�?             7@        ������������������������       �      �?              @        ������������������������       �                     .@        ������������������������       ��q�q�?             (@        �t�bh�h)h,K ��h.��R�(KKkKK��h\�B�       �{@     �p@     �v@     �U@     `u@     @U@               @     `u@     @S@     �t@     �Q@     0q@      D@     `m@      D@     �b@      ?@     �`@      7@     ``@      5@      F@      ,@     �U@      @     �S@      @      <@      @      ,@      �?      @              $@      �?      ,@      @     �I@      �?      B@              .@      �?       @       @      @       @      .@       @      @              "@       @     @U@      "@      D@      �?      .@      �?      @      �?       @              9@             �F@       @      B@       @      ,@       @      @       @       @              6@      @      @      @       @       @      @      �?      1@      @      @      �?      ,@       @       @              @       @      "@              D@             �M@      >@      @@      8@      5@      6@      4@      1@      1@      &@      @      @       @      @      @       @      (@      @      @      @      "@      �?      @      @      �?      @      &@       @      ;@      @      0@      @      @              "@      @      &@               @      @      9@       @      2@              @       @       @       @      @             @S@     �f@      @     @_@      @      D@              .@      @      9@       @      @      �?      2@              *@      �?      @             @U@     �R@      L@      "@      <@      @      @      @      7@              @      @      2@     @P@      <@     �A@      7@      <@      ,@      7@      @      3@      �?      &@               @      �?      @       @      @      &@      @      "@      @      @              @      >@      @      6@      �?      @      �?      .@               @      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ1�.hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsK}hth)h,K ��h.��R�(KK}��h{�B@         ,                 `f�$@�6��l�?�           @�@               !                    �?�iU��2�?�            0q@     "@                           �?9#��?�            @l@                                 �0@X�EQ]N�?�            �j@      @������������������������       �      �?              @                                  �;@�Q�1X�?�            �i@     @U@       
                   �9@�~t��?+            @Q@     D@       	                 �Y�@��a�n`�?'             O@      5@������������������������       ����Q��?             $@        ������������������������       � ��WV�?              J@      @������������������������       �և���X�?             @                                  �<@D��*�4�?U            @a@     T@                            @P�Lt�<�?-             S@      @������������������������       �                     (@      @                           �?      �?&             P@      @                        �Y�@      �?             @@       @������������������������       �                     (@Z      ������������������������       �ףp=
�?	             4@�      ������������������������       �                     @@�                                @@@��� ��?(             O@                               @3�@      �?             4@                              �?�@���|���?	             &@      ������������������������       �����X�?             @�      ������������������������       �      �?             @�      ������������������������       ������H�?             "@�                              �?�@@4և���?             E@      ������������������������       �                     7@                                @C@�S����?             3@       ������������������������       �                     @�      ������������������������       �      �?             (@(                                  8@"pc�
�?             &@       ������������������������       ��q�q�?             @J      ������������������������       �                     @3      "       +                    �?Tt�ó��?#            �H@      #       $                 ���@�G�z�?             D@        ������������������������       �@4և���?
             ,@�       %       (                    �?��
ц��?             :@        &       '                 �&B@�q�q�?	             "@       ������������������������       ����Q��?             @�       ������������������������       �      �?             @�       )       *                 �?�@��.k���?             1@        ������������������������       ��q�q�?             @�       ������������������������       ��eP*L��?             &@$       ������������������������       �                     "@       -       b                    �?��|���?           P{@       .       _                    @B.���?�            �o@       /       0                    $@�s�68e�?�            `l@        ������������������������       �                     1@�       1       V                    �?�������?�            @j@       2       A                     �?�ߥV��?m             e@        3       >                    �?�xGZ���?+            �Q@       4       =                   �L@X�<ݚ�?!             K@       5       <                 `f�B@�ݏ^���?            �F@       6       9                    ?@���Q��?             >@       7       8                   @>@���Q��?
             .@       ������������������������       ����!pc�?             &@`      ������������������������       �      �?             @:      :       ;                    G@z�G�z�?
             .@       ������������������������       ������H�?             "@?      ������������������������       ��q�q�?             @I      ������������������������       ��q�q�?             .@7      ������������������������       ������H�?             "@G       ?       @                    D@      �?
             0@      ������������������������       ��eP*L��?             &@!      ������������������������       ����Q��?             @�      B       O                   @<@ ���3�?B            �X@      C       H                 �R,@j�q����?&             I@        D       G                   �8@�q�q�?             .@      E       F                    5@z�G�z�?             $@       ������������������������       ����Q��?             @-      ������������������������       �                     @,      ������������������������       ����Q��?             @�      I       J                   �9@(N:!���?            �A@        ������������������������       �        
             *@�       K       N                    �?"pc�
�?             6@      L       M                 `fV7@���!pc�?	             &@      ������������������������       �z�G�z�?             @�      ������������������������       ��q�q�?             @�      ������������������������       ��C��2(�?             &@�      P       Q                 ���&@Hm_!'1�?            �H@       ������������������������       ��q�q�?             @�       R       U                    F@ �#�Ѵ�?            �E@      S       T                    D@�8��8��?             8@      ������������������������       ��}�+r��?             3@%      ������������������������       �z�G�z�?             @g      ������������������������       �                     3@�       W       \                   �B@������?            �D@       X       [                 �DpB@R���Q�?             4@       Y       Z                 �̌4@�8��8��?	             (@        ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ]       ^                   �J@���N8�?             5@       ������������������������       �                     *@        ������������������������       �      �?              @        `       a                    @ ��WV�?             :@        ������������������������       �؇���X�?             @        ������������������������       �                     3@        c       x                 �D�H@*
;&���?u             g@       d       w                    @��$�4��?K            �]@       e       l                     @�>4և��?F             \@       f       k                   �H@�U�=���?'            �P@       g       j                   �;@����˵�?"            �M@        h       i                    6@     ��?             @@        ������������������������       ����!pc�?             &@        ������������������������       �        	             5@        ������������������������       �                     ;@        ������������������������       �����X�?             @        m       v                    @�I� �?             G@       n       o                    @�θ�?            �C@        ������������������������       �                     *@        p       s                 ���0@$��m��?             :@       q       r                    �?������?             1@       ������������������������       ������H�?             "@        ������������������������       �      �?              @        t       u                    �?X�<ݚ�?             "@        ������������������������       ����Q��?             @        ������������������������       �      �?             @        ������������������������       �؇���X�?             @        ������������������������       �                     @        y       z                  "�b@Pa�	�?*            �P@       ������������������������       �                    �I@        {       |                    �?�r����?             .@       ������������������������       �                     $@        ������������������������       ����Q��?             @        �t�bh�h)h,K ��h.��R�(KK}KK��h\�B�       0{@     Pq@     �k@      K@     �h@      ;@     �g@      9@      @      @     `g@      4@     �M@      $@      L@      @      @      @      I@       @      @      @      `@      $@     �R@       @      (@              O@       @      >@       @      (@              2@       @      @@              K@       @      .@      @      @      @      @       @       @       @       @      �?     �C@      @      7@              0@      @      @              "@      @      "@       @      @       @      @              6@      ;@      *@      ;@      �?      *@      (@      ,@      @      @       @      @      �?      @      "@       @      @       @      @      @      "@             �j@     �k@     @g@     �P@      d@     �P@              1@      d@     �H@      _@     �F@      C@      @@      >@      8@      6@      7@      (@      2@      "@      @       @      @      �?      @      @      (@      �?       @       @      @      $@      @       @      �?       @       @      @      @      @       @     �U@      *@     �D@      "@      $@      @       @       @      @       @      @               @      @      ?@      @      *@              2@      @       @      @      @      �?      @       @      $@      �?     �F@      @      @       @     �D@       @      6@       @      2@      �?      @      �?      3@             �B@      @      1@      @      &@      �?      @      �?      @              @       @      4@      �?      *@              @      �?      9@      �?      @      �?      3@              <@     �c@      :@      W@      4@      W@      @     �N@      @      L@      @      =@      @       @              5@              ;@       @      @      .@      ?@      "@      >@              *@      "@      1@      @      *@      �?       @      @      @      @      @       @      @      @      �?      @      �?      @               @      P@             �I@       @      *@              $@       @      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJg�)hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKghth)h,K ��h.��R�(KKg��h{�B�         L                    �?<��z��?�           @�@                                  *@�>�S�?/           �~@       @                           @����"�?             =@      @������������������������       �                     2@      �?������������������������       �                     &@       @       1                   �<@8ӈ(�3�?            }@      @                           �?$s��O�?�            �q@      @                        ��.@�E��ӭ�?              K@      @	       
                    8@r�q��?             B@        ������������������������       �      �?             @     "@                        ��%@ףp=
�?             >@      @������������������������       �                     3@      7@������������������������       ����!pc�?             &@     �?                          �;@      �?             2@       ������������������������       ��n_Y�K�?             *@      @������������������������       �z�G�z�?             @       @                            �?�?v��?�            @l@                                 `@@������?             1@       ������������������������       ��q�q�?             @�      ������������������������       �                     &@w             &                   �;@X��J��?�             j@             %                    �?h��)�~�?D            @\@                              ���@���2j��?=            �Y@       ������������������������       �����X�?             ,@�             "                   �8@`���i��?6             V@                                  @P�2E��?*            @P@                                 �(@      �?             0@       ������������������������       �      �?              @      ������������������������       �                      @�                              @3�@@�E�x�?            �H@       ������������������������       �                     4@V              !                   �3@XB���?             =@       ������������������������       ������H�?             "@3      ������������������������       �                     4@A      #       $                     @�㙢�c�?             7@        ������������������������       �                     (@�       ������������������������       ����|���?             &@v       ������������������������       �                     &@j       '       0                    �? �q�q�?=             X@       (       /                 03�<@@�)�n�?6            @U@       )       *                     @�(\����?2             T@        ������������������������       ������H�?             "@�       +       ,                    �? ��PUp�?-            �Q@        ������������������������       �                     2@       -       .                 �?$@�O4R���?             �J@        ������������������������       ������H�?             "@-       ������������������������       �                     F@]       ������������������������       �z�G�z�?             @�       ������������������������       ��C��2(�?             &@A       2       ;                     �?
��^���?n            @g@        3       8                    �?�xGZ���?&            �Q@       4       5                    �?X�<ݚ�?            �F@        ������������������������       �      �?             (@�       6       7                 �T!@@4���C�?            �@@      ������������������������       ��q�q�?             8@�       ������������������������       �                     "@`      9       :                   �H@�q�����?             9@      ������������������������       �����X�?	             ,@;      ������������������������       �"pc�
�?             &@?      <       C                    @@�y��*�?H             ]@       =       @                    $@">�֕�?            �A@      >       ?                   �=@      �?             2@        ������������������������       ����Q��?             @      ������������������������       ���
ц��?             *@!      A       B                   �>@�t����?	             1@      ������������������������       �                      @�      ������������������������       ��<ݚ�?             "@8       D       K                   �*@ 7���B�?3            @T@      E       F                 �?�@ �h�7W�?$            �J@       ������������������������       �                     ;@-      G       J                    G@ȵHPS!�?             :@      H       I                 pFt @     ��?             0@       ������������������������       ��<ݚ�?             "@�       ������������������������       �؇���X�?             @�       ������������������������       �                     $@v      ������������������������       �                     <@�      M       b                   �=@���Y�?�             k@      N       Q                     @ XөM"�?]             a@       O       P                 ��*@�&=�w��?!            �J@       ������������������������       ��<ݚ�?             "@�      ������������������������       �                     F@�       R       a                 ��Y7@��6���?<             U@      S       ^                    �?և���X�?0            �O@      T       W                 ��@�eP*L��?#             F@       U       V                   @@�E��ӭ�?             2@       ������������������������       �؇���X�?             @�       ������������������������       ����|���?	             &@y       X       [                    �?
j*D>�?             :@       Y       Z                 �̌@      �?             0@        ������������������������       �      �?              @        ������������������������       �      �?              @        \       ]                   �9@�z�G��?
             $@        ������������������������       �z�G�z�?             @        ������������������������       ����Q��?             @        _       `                    �?p�ݯ��?             3@        ������������������������       �                      @        ������������������������       ����|���?             &@        ������������������������       ������?             5@        c       d                 `f$@      �?8             T@        ������������������������       ��q�q�?             @        e       f                     @�L���?3            �R@       ������������������������       �        -            �P@        ������������������������       �      �?              @        �t�bh�h)h,K ��h.��R�(KKgKK��h\�Bp       p|@     p@     �x@     �X@      &@      2@              2@      &@              x@      T@     �n@      A@     �C@      .@      >@      @      @      @      ;@      @      3@               @      @      "@      "@      @       @      @      �?     �i@      3@      *@      @       @      @      &@             @h@      .@     �Y@      &@     �V@      &@      $@      @     @T@      @      O@      @      ,@       @      @       @       @              H@      �?      4@              <@      �?       @      �?      4@              3@      @      (@              @      @      &@              W@      @     �T@      @     �S@       @       @      �?     �Q@      �?      2@              J@      �?       @      �?      F@              @      �?      $@      �?     �a@      G@      C@      @@      9@      4@      @      @      3@      ,@      $@      ,@      "@              *@      (@      @      $@      "@       @     �Y@      ,@      8@      &@      "@      "@       @      @      @      @      .@       @       @              @       @     �S@      @      I@      @      ;@              7@      @      *@      @      @       @      @      �?      $@              <@              M@     �c@      H@     @V@       @     �I@       @      @              F@      G@      C@      ;@      B@      4@      8@      @      *@      �?      @      @      @      .@      &@      (@      @      @      @      @      �?      @      @      �?      @       @      @      @      (@               @      @      @      3@       @      $@     �Q@      @       @      @      Q@             �P@      @       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�]_AhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKkhth)h,K ��h.��R�(KKk��h{�B�         Z                  x#J@~�Я��?�           @�@              9                    �?j;v�>��?x           ��@    �@@                        ���"@�#߆;s�?            z@                                    @�?�<��?�            `h@      �?������������������������       �                     &@                                   �?�LQ�1	�?x             g@     @                          �;@󝢸]�?q            �e@       @                          �7@d��0u��?%             N@     �?	       
                   �5@��r._�?            �D@       ������������������������       ���a�n`�?             ?@      @������������������������       �                     $@                                  �8@�����?             3@      T@������������������������       ����Q��?             $@      @������������������������       ��<ݚ�?             "@      @                          �<@x�}b~|�?L            �\@      @                        �?�@�O4R���?$            �J@      @������������������������       �                     E@Z      ������������������������       ��C��2(�?             &@�                                 �?f>�cQ�?(            �N@                                 @@@�t����?             1@       ������������������������       �����X�?             @n      ������������������������       �                     $@�      ������������������������       ��C��2(�?             F@�      ������������������������       �ףp=
�?             $@�                                 *@$~���?�            �k@                                  @4���C�?            �@@      ������������������������       �                     0@                              ��T?@@�0�!��?
             1@      ������������������������       �                      @�      ������������������������       ��q�q�?             "@(             8                    �?�S����?o            �g@              #                   �9@Ld����?[            �c@       !       "                   �3@`2U0*��?             9@       ������������������������       �r�q��?             @A      ������������������������       �                     3@�       $       5                   �>@��T�l��?K            �`@       %       4                 ���=@"��$�?@            �[@       &       -                   �=@�����?:            �X@        '       *                 ��\,@<=�,S��?            �A@        (       )                   �'@��
ц��?             *@        ������������������������       �և���X�?             @�       ������������������������       ��q�q�?             @�       +       ,                    �?���!pc�?             6@        ������������������������       ����Q��?             $@       ������������������������       �r�q��?             (@       .       1                   �I@�����H�?$            �O@       /       0                 ��$:@�MI8d�?            �B@       ������������������������       �h�����?             <@�       ������������������������       �X�<ݚ�?             "@A       2       3                   �N@ ��WV�?             :@       ������������������������       �                     3@�       ������������������������       �؇���X�?             @�       ������������������������       ��n_Y�K�?             *@�       6       7                   �C@���N8�?             5@      ������������������������       �                     ,@�       ������������������������       �؇���X�?             @`      ������������������������       �                    �@@:      :       W                    @b����?t            �g@      ;       F                 `f�%@�q�q�?l             e@       <       C                 pF @�>���?%             K@      =       @                    �?�������?             A@      >       ?                 ���@��<b���?             7@        ������������������������       �      �?              @      ������������������������       ���S�ۿ?
             .@!      A       B                    8@���|���?             &@       ������������������������       �����X�?             @�      ������������������������       �      �?             @8       D       E                   �5@z�G�z�?             4@       ������������������������       �և���X�?             @      ������������������������       �$�q-�?	             *@-      G       N                     @���y4F�?G            �\@      H       I                     �?г�wY;�?+             Q@       ������������������������       ������H�?             "@�       J       M                   �*@P����?%            �M@        K       L                    =@�X�<ݺ?             2@      ������������������������       ������H�?             "@�      ������������������������       �                     "@�      ������������������������       �                    �D@�      O       R                    �?
;&����?             G@       P       Q                 ��.@     ��?             0@       ������������������������       �X�<ݚ�?             "@�       ������������������������       �                     @      S       V                 ���4@*;L]n�?             >@      T       U                    �?�����?             3@       ������������������������       �X�<ݚ�?             "@g      ������������������������       �ףp=
�?             $@�       ������������������������       �                     &@y       X       Y                   �0@��s����?             5@        ������������������������       �                     &@�       ������������������������       ����Q��?             $@        [       h                    �?lwY���?B            @Z@       \       c                    �?r�q��?6             U@        ]       b                    �?���|���?            �@@       ^       _                   �;@և���X�?             5@        ������������������������       ��<ݚ�?             "@        `       a                  �}S@�q�q�?             (@        ������������������������       �      �?             @        ������������������������       ��q�q�?             @        ������������������������       �      �?             (@        d       g                   �:@`'�J�?!            �I@        e       f                    �?z�G�z�?	             $@       ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                    �D@        i       j                    :@؇���X�?             5@        ������������������������       ����Q��?             @        ������������������������       �                     0@        �t�bh�h)h,K ��h.��R�(KKkKK��h\�B�       �{@     �p@     �y@     �h@     �u@     @R@     `e@      8@      &@              d@      8@     �b@      7@     �G@      *@      A@      @      8@      @      $@              *@      @      @      @      @       @      Z@      $@      J@      �?      E@              $@      �?      J@      "@      (@      @       @      @      $@              D@      @      "@      �?     �e@     �H@      ,@      3@              0@      ,@      @       @              @      @      d@      >@     �_@      >@      8@      �?      @      �?      3@             �Y@      =@     �T@      <@     �S@      4@      6@      *@      @      @      @      @       @      @      0@      @      @      @      $@       @      L@      @      ?@      @      ;@      �?      @      @      9@      �?      3@              @      �?      @       @      4@      �?      ,@              @      �?     �@@             �P@     �^@     �H@     �]@      9@      =@      "@      9@      @      2@      @      @      �?      ,@      @      @       @      @       @       @      0@      @      @      @      (@      �?      8@     �V@       @     �P@      �?       @      �?      M@      �?      1@      �?       @              "@             �D@      6@      8@      @      &@      @      @              @      1@      *@      @      *@      @      @      �?      "@      &@              1@      @      &@              @      @      @@     @R@      ,@     �Q@      (@      5@      "@      (@       @      @      @      @      @      @      @       @      @      "@       @     �H@       @       @              @       @       @             �D@      2@      @       @      @      0@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJL�OhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsK{hth)h,K ��h.��R�(KK{��h{�B�         d                  x#J@������?�           @�@                                  @,˫�5�?�           ��@ �3	�                             @��a�n`�?             ?@       ������������������������       �                     3@        ������������������������       ��q�q�?             (@      @       5                  �#@� :N?��?o           ��@      �?                           /@6�	�j��?�            `q@      @������������������������       �z�G�z�?             @      >@	       4                    �?��0%�?�            q@       
       %                   �<@tMI!>�?�            �k@     "@       "                    �?��a�n`�?a            `c@      @                          �;@dP-���?Y            �a@     7@                        ��Y@������?.            �Q@      �?������������������������       ��q�q�?             @                                 �0@     p�?*             P@      @������������������������       �z�G�z�?             $@       @                        �?$@�X�<ݺ?&             K@       ������������������������       �        
             *@�                              �{@��p\�?            �D@       ������������������������       �r�q��?             @w                              @3�@ >�֕�?            �A@       ������������������������       �        	             (@�                                �3@���}<S�?             7@       ������������������������       �r�q��?             @�      ������������������������       ��IєX�?
             1@�             !                 �?$@0z�(>��?+            �Q@                                  @�L���?            �B@       ������������������������       �                     @                                  �?��a�n`�?             ?@                              ���@HP�s��?             9@      ������������������������       �      �?             0@V      ������������������������       �                     "@J      ������������������������       �r�q��?             @3      ������������������������       �                     A@A      #       $                   �9@d}h���?             ,@        ������������������������       �      �?             @�       ������������������������       �                      @v       &       )                    �?@�0�!��?,             Q@        '       (                    @@     ��?             0@        ������������������������       ����Q��?             @�       ������������������������       �                     &@�       *       +                 �&B@D>�Q�?!             J@        ������������������������       �                     .@$       ,       1                 ��i @���"͏�?            �B@       -       .                 �?�@�	j*D�?             :@        ������������������������       �r�q��?             (@-       /       0                   �@@և���X�?	             ,@       ������������������������       �      �?             @�       ������������������������       �      �?              @A       2       3                   �A@�C��2(�?             &@        ������������������������       �r�q��?             @�       ������������������������       �                     @�       ������������������������       ����Q��?             I@�       6       Q                    �?l~X���?�             r@      7       P                   �K@�q�qT�?|             h@       8       ;                    ,@�ݿ���?s            `f@       9       :                    �?ҳ�wY;�?
             1@       ������������������������       �r�q��?             @;      ������������������������       ��eP*L��?             &@?      <       G                 ��D:@�$�����?i            @d@      =       >                    �?�8��8��?D             [@       ������������������������       ����|���?	             &@G       ?       @                   �;@h�a��?;            @X@       ������������������������       �                    �B@!      A       D                   @@@�8��8��?$             N@       B       C                    �?r�q��?             2@       ������������������������       �؇���X�?             @8       ������������������������       �"pc�
�?             &@8      E       F                   �*@���N8�?             E@       ������������������������       ��<ݚ�?             "@-      ������������������������       �                    �@@,      H       O                    �?�{��?��?%             K@      I       L                   �>@�5��
J�?              G@       J       K                 ��=@��}*_��?             ;@        ������������������������       �z�G�z�?	             .@v      ������������������������       ��q�q�?	             (@�      M       N                 `f�B@�}�+r��?             3@       ������������������������       �r�q��?             @�      ������������������������       �        
             *@�      ������������������������       �                      @�      ������������������������       ��n_Y�K�?	             *@�       R       U                   �0@�q�q��?E             X@       S       T                 `f�=@�8��8��?             (@       ������������������������       �      �?             @%      ������������������������       �                      @g      V       ]                     @d}h���?=             U@       W       Z                    6@,�+�C�?)            �K@        X       Y                   �;@�����H�?             ;@        ������������������������       ��θ�?	             *@�       ������������������������       �                     ,@        [       \                   �H@h�����?             <@       ������������������������       �                     7@        ������������������������       �z�G�z�?             @        ^       c                 `v�6@l��[B��?             =@       _       b                 03�1@�X����?             6@       `       a                 ��.@      �?             0@        ������������������������       ����Q��?             @        ������������������������       �"pc�
�?             &@        ������������������������       �      �?             @        ������������������������       �                     @        e       x                     �?84(���?I            �\@       f       q                    �?r٣����??            �X@        g       n                    �?8����?             G@       h       m                   @E@     ��?             @@       i       j                 ��+T@���y4F�?             3@        ������������������������       �                     @        k       l                    =@�	j*D�?             *@       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       ��n_Y�K�?             *@        o       p                   �D@X�Cc�?             ,@        ������������������������       �؇���X�?             @        ������������������������       �և���X�?             @        r       u                    �?r�����?!            �J@        s       t                    �?���Q��?             .@       ������������������������       ��eP*L��?             &@        ������������������������       �      �?             @        v       w                    �?P�Lt�<�?             C@       ������������������������       �                     @@        ������������������������       �r�q��?             @        y       z                    �?      �?
             0@        ������������������������       ����|���?             &@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK{KK��h\�B�        |@     `p@     �y@     �f@      @      8@              3@      @      @     py@     �c@      k@     �N@      �?      @      k@     �L@     �h@      ;@     �a@      .@      `@      (@     �N@      "@       @      @     �M@      @       @       @     �I@      @      *@              C@      @      @      �?     �@@       @      (@              5@       @      @      �?      0@      �?      Q@      @      A@      @      @              <@      @      7@       @      ,@       @      "@              @      �?      A@              &@      @      @      @       @              L@      (@      *@      @       @      @      &@             �E@      "@      .@              <@      "@      2@       @      $@       @       @      @      @      @      @      @      $@      �?      @      �?      @              4@      >@     �g@     �X@      d@      ?@      c@      :@      &@      @      @      �?      @      @     �a@      4@     �X@      "@      @      @      W@      @     �B@             �K@      @      .@      @      @      �?      "@       @      D@       @      @       @     �@@             �E@      &@     �A@      &@      1@      $@      (@      @      @      @      2@      �?      @      �?      *@               @               @      @      =@     �P@      &@      �?      @      �?       @              2@     �P@      @     �I@      @      8@      @      $@              ,@      �?      ;@              7@      �?      @      ,@      .@      @      .@      @      (@       @      @       @      "@      @      @      @              B@     �S@      8@     �R@      ,@      @@      "@      7@      @      .@              @      @      "@      @      @              @      @       @      @      "@      �?      @      @      @      $@     �E@      "@      @      @      @      @      �?      �?     �B@              @@      �?      @      (@      @      @      @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ��lhG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKohth)h,K ��h.��R�(KKo��h{�B�         (                     @4�<����?�           @�@                                   �?x����?�            �r@                                  (@x���@O�?o             e@        ������������������������       �                     "@                                   �?��Q���?h             d@      �?                        pVAH@<ݚ)�?             B@     �?       
                    �?z�G�z�?             9@              	                 ���<@�t����?             1@        ������������������������       ��<ݚ�?             "@       ������������������������       �      �?              @      @������������������������       �                      @                                  �8@�eP*L��?             &@      T@������������������������       �      �?             @      @������������������������       �����X�?             @      @                          @>@���-T��?P             _@     @                           &@XI�~�?2            @S@       @������������������������       �      �?             0@Z                              ��D:@�.ߴ#�?&            �N@                                �*@�(\����?             D@       ������������������������       ��}�+r��?             3@w      ������������������������       �                     5@n                                 J@�����?             5@      ������������������������       �r�q��?             (@�      ������������������������       �                     "@�                                 @@�7����?            �G@       ������������������������       �r�q��?             @c      ������������������������       �� ��1�?            �D@             #                   �;@���f�?Y             `@                                   �?�:�]��?!            �I@                                 6@�X�<ݺ?             B@       ������������������������       �"pc�
�?             &@V      ������������������������       �                     9@J      !       "                 ��J@�r����?             .@      ������������������������       �                     $@A      ������������������������       ����Q��?             @�       $       '                     �?�(�Tw�?8            �S@       %       &                 0��I@P�Lt�<�?             C@        ������������������������       �      �?             @j       ������������������������       �                     A@�       ������������������������       �                     D@�       )       n                    @�G�5��?�            �y@       *       +                    �?.��<�?�             y@        ������������������������       �؇���X�?             ,@$       ,       U                    �?���0���?�            @x@       -       2                   �0@$G$n��?�            0p@        .       /                    !@ҳ�wY;�?             A@        ������������������������       ��E��ӭ�?             2@]       0       1                    *@     ��?             0@        ������������������������       ����Q��?             @A       ������������������������       ����|���?             &@�       3       <                  ��@�W�l~�?�             l@        4       ;                 �Y�@�i�y�?+            �O@       5       :                 ���@�7��?            �C@       6       7                    �?(;L]n�?             >@       ������������������������       �                     $@�       8       9                 ��@P���Q�?             4@      ������������������������       ��C��2(�?             &@:      ������������������������       �                     "@;      ������������������������       ������H�?             "@?      ������������������������       �                     8@I      =       @                   @@H�ՠ&��?h            @d@       >       ?                 �?$@����X�?             5@       ������������������������       �      �?             0@      ������������������������       ����Q��?             @!      A       N                   �<@�*/�8V�?X            �a@      B       C                 �?�@�7��d��?>             Y@       ������������������������       �                    �A@8       D       I                 ���!@ ����?)            @P@       E       H                   �;@r�q��?             >@      F       G                 ��Y @����X�?
             ,@       ������������������������       ����Q��?             @,      ������������������������       ��<ݚ�?             "@�      ������������������������       �      �?	             0@�       J       M                    ;@ >�֕�?            �A@        K       L                 ��q1@z�G�z�?             $@       ������������������������       �                     @�      ������������������������       ����Q��?             @�      ������������������������       �                     9@�      O       R                   @@@� ��1�?            �D@       P       Q                    ?@�q�q�?             (@       ������������������������       �և���X�?             @�       ������������������������       �z�G�z�?             @      S       T                   �D@XB���?             =@      ������������������������       �                     8@%      ������������������������       �z�G�z�?             @g      V       ]                    �?&X�IN�?K             `@        W       X                    �?�q�q�?            �C@        ������������������������       �և���X�?             @}       Y       Z                    9@     ��?             @@        ������������������������       �z�G�z�?             $@        [       \                 �&B@�X����?             6@       ������������������������       �X�Cc�?	             ,@        ������������������������       �      �?              @        ^       k                 ���4@$�ݏ^��?3            �V@       _       j                   @B@`՟�G��?$             O@       `       i                    �?      �?              L@       a       f                 ��&@(옄��?             G@       b       e                 @3�@�c�Α�?             =@       c       d                 �&B@b�2�tk�?
             2@        ������������������������       �և���X�?             @        ������������������������       ����|���?             &@        ������������������������       ��C��2(�?             &@        g       h                    =@������?             1@        ������������������������       �����X�?             @        ������������������������       �z�G�z�?             $@        ������������������������       ��z�G��?             $@        ������������������������       �                     @        l       m                    !@h�����?             <@        ������������������������       �r�q��?             @        ������������������������       �                     6@        ������������������������       �                     (@        �t�bh�h)h,K ��h.��R�(KKoKK��h\�B�        |@     �p@      a@     @d@     ``@      C@              "@     ``@      =@      9@      &@      4@      @      (@      @      @       @      @      @       @              @      @      @      �?       @      @     �Z@      2@      R@      @      ,@       @      M@      @     �C@      �?      2@      �?      5@              3@       @      $@       @      "@              A@      *@      �?      @     �@@       @      @      _@      @     �G@       @      A@       @      "@              9@       @      *@              $@       @      @      �?     @S@      �?     �B@      �?      @              A@              D@     �s@     �Y@     �r@     �Y@       @      (@     �r@     �V@      l@     �A@      6@      (@      *@      @      "@      @       @      @      @      @     @i@      7@     �N@       @     �B@       @      =@      �?      $@              3@      �?      $@      �?      "@               @      �?      8@             �a@      5@      .@      @      (@      @      @       @     �_@      .@     @W@      @     �A@              M@      @      9@      @      $@      @      @       @      @       @      .@      �?     �@@       @       @       @      @              @       @      9@             �@@       @      @      @      @      @      �?      @      <@      �?      8@              @      �?     �R@     �K@      *@      :@      @      @      "@      7@       @       @      @      .@      @      "@       @      @     �N@      =@      A@      <@      <@      <@      9@      5@      5@       @      &@      @      @      @      @      @      $@      �?      @      *@       @      @       @       @      @      @      @              ;@      �?      @      �?      6@              (@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�-#hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKwhth)h,K ��h.��R�(KKw��h{�B�         R                    �?4�<����?�           @�@                                  @$�|:	�?%           �~@                                    @����X�?             <@       ������������������������       �        
             3@        ������������������������       ������H�?             "@      �?       ;                 ��i=@z�#��o�?           �|@                               �1@`�3Ka��?�            �u@      _@                          �;@��H�??             W@      9@	                          �8@h+�v:�?             A@       
                           �?��<b���?             7@      "@������������������������       �      �?              @      @������������������������       �                     .@     7@������������������������       ����!pc�?             &@      �?                           �? 	��p�?(             M@                                ���@PN��T'�?             ;@      @������������������������       �                     @       @������������������������       ���s����?             5@Z      ������������������������       �                     ?@�             8                    �?�"$����?�            0p@                                 �?(.��H�?�            `m@                                 �<@XB���?             =@                                  @P���Q�?             4@       ������������������������       �r�q��?             @�      ������������������������       �        	             ,@�      ������������������������       �                     "@�             5                    �?8�Jh�a�?x            �i@             (                     @���'\�?j            �f@                               `f�)@"pc�
�?"            �K@                                  =@@4և���?	             ,@       ������������������������       �؇���X�?             @(      ������������������������       �                     @V              %                 ��$:@��P���?            �D@      !       $                   �*@�+$�jP�?             ;@      "       #                   �;@�d�����?             3@       ������������������������       �                     $@�       ������������������������       �X�<ݚ�?             "@�       ������������������������       �                      @v       &       '                   `G@����X�?             ,@        ������������������������       ������H�?             "@�       ������������������������       ����Q��?             @�       )       0                    ?@�m(']�?H            �_@       *       +                 @3�@�|���?5             V@        ������������������������       �                    �@@$       ,       /                 ��Y @ �Jj�G�?             �K@       -       .                   �5@�nkK�?             7@        ������������������������       �z�G�z�?             @-       ������������������������       �                     2@]       ������������������������       �                     @@�       1       2                   @@@��-�=��?            �C@        ������������������������       ��<ݚ�?             "@�       3       4                 @3�@��S�ۿ?             >@        ������������������������       �8�Z$���?             *@�       ������������������������       �                     1@�       6       7                    >@�8��8��?             8@      ������������������������       �                     ,@�       ������������������������       �z�G�z�?             $@`      9       :                    0@�q�q�?             8@       ������������������������       �X�<ݚ�?             "@;      ������������������������       �                     .@?      <       K                    �?�X����?=            �[@      =       @                   �>@rr�J��?(            �R@       >       ?                   �<@`�Q��?
             9@        ������������������������       �                     (@      ������������������������       ��n_Y�K�?             *@!      A       D                    �? \� ���?            �H@       B       C                  �}S@      �?
             0@       ������������������������       �z�G�z�?             @8       ������������������������       ����|���?             &@8      E       J                 03S@<���D�?            �@@      F       I                   �B@`2U0*��?             9@      G       H                    �?�C��2(�?
             &@      ������������������������       �r�q��?             @�      ������������������������       �                     @�       ������������������������       �                     ,@�       ������������������������       �      �?              @v      L       O                 ��H@r�q��?             B@      M       N                     @���N8�?             5@      ������������������������       �@4և���?             ,@�      ������������������������       �                     @�      P       Q                    �?�q�q�?
             .@      ������������������������       �z�G�z�?             $@�       ������������������������       ����Q��?             @      S       b                     @� �th}�?�            �k@      T       _                  "�b@`Jj��?M             _@      U       Z                    �?����?B            �Z@       V       Y                     �? �Cc}�?             <@       W       X                   �H@�S����?             3@       ������������������������       �                     *@}       ������������������������       �      �?             @�       ������������������������       �                     "@        [       ^                   �;@ ���J��?1            �S@        \       ]                    6@�C��2(�?             6@        ������������������������       ����Q��?             @        ������������������������       �                     1@        ������������������������       �                      L@        `       a                    <@r�q��?             2@        ������������������������       ��q�q�?             "@        ������������������������       �                     "@        c       r                   �<@�fSO��?E            �X@       d       o                    @F~��7�?9            �T@       e       j                    �?ޚ)�?1             R@       f       g                 ��@���j��?!             G@        ������������������������       �ףp=
�?             4@        h       i                    �?
j*D>�?             :@       ������������������������       �D�n�3�?             3@        ������������������������       �                     @        k       l                 pF�-@��
ц��?             :@        ������������������������       �                      @        m       n                 ��1@�<ݚ�?             2@        ������������������������       �                     "@        ������������������������       �X�<ݚ�?             "@        p       q                  �:@�C��2(�?             &@        ������������������������       �z�G�z�?             @        ������������������������       �                     @        s       t                   �>@     ��?             0@        ������������������������       �      �?              @        u       v                    �?      �?              @        ������������������������       �      �?             @        ������������������������       �      �?             @        �t�b���      h�h)h,K ��h.��R�(KKwKK��h\�Bp        |@     �p@     �x@     �W@       @      4@              3@       @      �?      x@     �R@     ps@      D@     �R@      1@      5@      *@      2@      @      @      @      .@              @       @      K@      @      7@      @      @              1@      @      ?@             �m@      7@      k@      2@      <@      �?      3@      �?      @      �?      ,@              "@             �g@      1@     �d@      .@     �F@      $@      *@      �?      @      �?      @              @@      "@      6@      @      ,@      @      $@              @      @       @              $@      @       @      �?       @      @     �^@      @     �U@      �?     �@@              K@      �?      6@      �?      @      �?      2@              @@             �A@      @      @       @      <@       @      &@       @      1@              6@       @      ,@               @       @      3@      @      @      @      .@             �R@     �A@     �F@      =@       @      1@              (@       @      @     �B@      (@       @       @      �?      @      @      @      =@      @      8@      �?      $@      �?      @      �?      @              ,@              @      @      >@      @      4@      �?      *@      �?      @              $@      @       @       @       @      @      K@      e@       @      ]@      @     @Y@      @      9@      @      0@              *@      @      @              "@       @      S@       @      4@       @      @              1@              L@      @      .@      @      @              "@      G@     �J@     �A@      H@      9@     �G@      *@     �@@       @      2@      &@      .@      &@       @              @      (@      ,@       @              @      ,@              "@      @      @      $@      �?      @      �?      @              &@      @      @      �?      @      @       @       @       @       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ5�;5hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsK_hth)h,K ��h.��R�(KK_��h{�B�                             @@cF �?�           @�@                                03�:@�p ��?            �D@                               ��k'@ �q�q�?             8@        ������������������������       �      �?              @      @������������������������       �                     0@      2@                           @�t����?             1@        ������������������������       ��C��2(�?             &@      $@������������������������       ��q�q�?             @      "@	       D                    �?TK;����?�           ��@       
       A                 Ј�U@��u�T(�?(           p|@     @                            �?��r>�?           `{@                                  �E@h��Q(�?/            �P@     T@                          �;@*O���?             B@      @������������������������       �      �?             @      @                          �B@     ��?             @@     @                          @>@�eP*L��?             6@      @������������������������       �     ��?             0@Z      ������������������������       �r�q��?             @�      ������������������������       �                     $@�                              �UwR@�g�y��?             ?@      ������������������������       �                     7@n      ������������������������       �      �?              @�                                  @ c�^��?�            0w@                                  �?����?�?;            �V@                              `fF)@      �?*             P@       ������������������������       �                     9@c      ������������������������       ��7��?            �C@      ������������������������       �                     :@             *                    �?h?\P��?�            �q@              !                   �7@D��\��?,            �Q@                                  �3@���|���?
             &@      ������������������������       �؇���X�?             @J      ������������������������       �      �?             @3      "       #                  ��@ףp=
�?"             N@       ������������������������       �                     >@�       $       )                    �?z�G�z�?             >@       %       (                    >@      �?             8@       &       '                 ��(@�����?             3@        ������������������������       ����|���?             &@�       ������������������������       �      �?              @�       ������������������������       �                     @�       ������������������������       �                     @�       +       ,                   `@��S�ۿ?�            @j@        ������������������������       �      �?              @       -       @                 �T�I@(a��䛼?�            @i@       .       7                   �<@h�a��?            @h@       /       0                   �0@�ㄡ^�?X             a@        ������������������������       ��8��8��?             (@�       1       4                   �:@��v��?P            @_@       2       3                 �1@ ��PUp�?.            �Q@        ������������������������       � 7���B�?             ;@�       ������������������������       �                     F@�       5       6                    �? 7���B�?"             K@       ������������������������       �`Ӹ����?            �F@      ������������������������       �                     "@�       8       ;                   @@@�KM�]�?'            �L@       9       :                   �>@X�Cc�?
             ,@       ������������������������       �؇���X�?             @;      ������������������������       �և���X�?             @?      <       =                   �E@ qP��B�?            �E@      ������������������������       �                     <@7      >       ?                    G@��S�ۿ?
             .@        ������������������������       �z�G�z�?             @      ������������������������       �                     $@!      ������������������������       �      �?              @�      B       C                    �?��.k���?
             1@       ������������������������       �؇���X�?             @8       ������������������������       ��z�G��?             $@8      E       T                 `f�%@����|e�?�             k@       F       I                 ���@     8�?)             P@       G       H                 03s@�����?	             5@       ������������������������       �z�G�z�?             @�      ������������������������       �      �?             0@�       J       K                    �?�K��&�?             �E@        ������������������������       ��n_Y�K�?             *@v      L       O                 `�X!@�q�q�?             >@       M       N                   �6@������?             .@       ������������������������       �      �?             @�      ������������������������       ������H�?             "@�      P       S                    �?���Q��?             .@      Q       R                   �:@���Q��?             $@        ������������������������       ����Q��?             @      ������������������������       �z�G�z�?             @-      ������������������������       �                     @%      U       X                     @��.��?^             c@      V       W                 ���a@�?�|�?C            �[@       ������������������������       �        <             Y@y       ������������������������       ����!pc�?             &@}       Y       ^                    �?D^��#��?            �D@       Z       [                    �?�q�q�?             ;@        ������������������������       �8�Z$���?             *@        \       ]                 ��*4@      �?             ,@        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �@4և���?             ,@        �t�bh�h)h,K ��h.��R�(KK_KK��h\�B�       }@     �n@      @     �A@      �?      7@      �?      @              0@      @      (@      �?      $@      @       @     �|@     �j@     py@      H@     �x@      D@     �J@      ,@      7@      *@      �?      @      6@      $@      (@      $@      &@      @      �?      @      $@              >@      �?      7@              @      �?     �u@      :@      V@       @      O@       @      9@             �B@       @      :@             p@      8@     �N@      $@      @      @      @      �?      �?      @      K@      @      >@              8@      @      2@      @      *@      @      @      @      @       @      @              @             �h@      ,@      @       @     �g@      (@      g@      $@     �`@      @      &@      �?     �^@      @     �Q@      �?      :@      �?      F@              J@       @     �E@       @      "@             �I@      @      "@      @      @      �?      @      @      E@      �?      <@              ,@      �?      @      �?      $@              @       @      "@       @      @      �?      @      @      J@     �d@      ;@     �B@       @      3@      �?      @      �?      .@      9@      2@      @       @      4@      $@      &@      @      @      @       @      �?      "@      @      @      @      @       @      �?      @      @              9@     �_@      @      [@              Y@      @       @      6@      3@      "@      2@       @      &@      @      @      �?      @      @              *@      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJi4�hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKmhth)h,K ��h.��R�(KKm��h{�B@         2                     @�)�>_M�?�           @�@               %                    �?0�矆��?�            �t@                                  �?j�'�=z�?~            �h@                               ��$:@�9���[�?S            �_@     �?                        `f�)@���Ls�?,            @P@      �?������������������������       �                     9@       @                          �;@R���Q�?             D@        ������������������������       �                     &@      �?	                        ���+@V�a�� �?             =@       
                          @B@�q�q�?             2@       ������������������������       ����|���?             &@        ������������������������       �����X�?             @        ������������������������       �                     &@                                �U�R@�ɞ`s�?'            �N@                               �DHC@t�F�}�?!            �I@                                  D@��Q��?             D@                                 �<@
;&����?             7@                                  �?և���X�?
             ,@        ������������������������       ����Q��?             @        ������������������������       �X�<ݚ�?             "@        ������������������������       �X�<ݚ�?             "@        ������������������������       ��t����?             1@        ������������������������       �                     &@        ������������������������       �      �?             $@                                   :@*O���?+             R@                                   9@D�n�3�?             3@        ������������������������       �և���X�?             @        ������������������������       ��q�q�?             (@               $                    �?�#ʆA��?            �J@                                 �;@���N8�?             E@        ������������������������       �      �?              @                !                   @B@�t����?             A@        ������������������������       �                     *@3      "       #                   @H@��s����?             5@      ������������������������       ����Q��?             $@�       ������������������������       �                     &@�       ������������������������       ��eP*L��?             &@v       &       /                    �?��ɉ�?U            @`@       '       .                    �?@�)�n�?:            @U@       (       +                     �? �h�7W�?%            �J@       )       *                    G@ 7���B�?             ;@       ������������������������       �                     7@�       ������������������������       �      �?             @$       ,       -                    =@$�q-�?             :@        ������������������������       �z�G�z�?             $@       ������������������������       �                     0@-       ������������������������       �                     @@]       0       1                     �?����?�?            �F@        ������������������������       ��IєX�?
             1@A       ������������������������       �                     <@�       3       X                    �?�q�q*�?�             x@       4       W                 �T�I@0Lj����?�             q@       5       R                   @@@���B��?�            pp@       6       7                    �?,���α�?�            �j@       ������������������������       �f���M�?             ?@�       8       O                   �<@L�)>|�?q            �f@      9       N                    �?����q �?b             d@      :       M                    0@�d�g��?W            �a@      ;       >                    �?|�(��?O            �_@       <       =                  ��@�X�<ݺ?             2@       ������������������������       �                     @7      ������������������������       ��8��8��?             (@G       ?       @                   �0@�����H�?D             [@       ������������������������       �����X�?             @!      A       B                   �3@�L�L��??            @Y@       ������������������������       �        
             7@�      C       D                   �4@�:�^���?5            �S@        ������������������������       ��q�q�?             @8      E       H                 �1@�n���?0             R@       F       G                 ��@���y4F�?             3@      ������������������������       �$�q-�?             *@,      ������������������������       �      �?             @�      I       J                 ��) @�O4R���?$            �J@       ������������������������       �                    �C@�       K       L                    :@@4և���?
             ,@       ������������������������       �                     @�      ������������������������       ������H�?             "@�      ������������������������       �                     ,@�      ������������������������       �                     5@�      P       Q                 @3�@8�A�0��?             6@      ������������������������       ���
ц��?             *@�       ������������������������       ��<ݚ�?             "@      S       T                 �?�@@�E�x�?"            �H@      ������������������������       �                     <@%      U       V                 pF� @���N8�?             5@       ������������������������       �      �?              @�       ������������������������       �        	             *@y       ������������������������       �X�<ݚ�?             "@}       Y       l                 `v�6@�Cc}��?K             \@       Z       g                    �?���!���??            �W@       [       d                    �?\X��t�?-            @Q@       \       _                    �?Fx$(�?             I@       ]       ^                    9@      �?             <@        ������������������������       �                      @        ������������������������       ���Q��?             4@        `       a                 ��@�eP*L��?             6@        ������������������������       ����Q��?             @        b       c                   �9@j���� �?             1@        ������������������������       �                     "@        ������������������������       �      �?              @        e       f                    .@D�n�3�?             3@        ������������������������       �                     "@        ������������������������       �z�G�z�?             $@        h       i                 ���.@z�G�z�?             9@        ������������������������       ��q�q�?	             (@        j       k                 03c4@$�q-�?	             *@       ������������������������       �                     @        ������������������������       �r�q��?             @        ������������������������       �                     2@        �t�bh�h)h,K ��h.��R�(KKmKK��h\�B�       `{@      q@     �b@      f@     `b@     �I@     @Y@      9@     �M@      @      9@              A@      @      &@              7@      @      (@      @      @      @      @       @      &@              E@      3@     �B@      ,@      :@      ,@      &@      (@      @       @       @      @      @      @      @      @      .@       @      &@              @      @      G@      :@       @      &@      @      @      @       @      C@      .@      @@      $@       @      @      >@      @      *@              1@      @      @      @      &@              @      @      @     �_@      @     �T@      @      I@      �?      :@              7@      �?      @       @      8@       @       @              0@              @@      �?      F@      �?      0@              <@     �q@     @X@     @m@      C@     �l@      A@     �f@     �@@      4@      &@      d@      6@     �b@      *@     �_@      *@     @\@      *@      1@      �?      @              &@      �?      X@      (@       @      @     �W@      @      7@             �Q@      @      @       @     �P@      @      .@      @      (@      �?      @      @      J@      �?     �C@              *@      �?      @               @      �?      ,@              5@              *@      "@      @      @      @       @      H@      �?      <@              4@      �?      @      �?      *@              @      @     �J@     �M@     �A@     �M@      >@     �C@      3@      ?@      @      5@               @      @      *@      (@      $@       @      @      $@      @      "@              �?      @      &@       @      "@               @       @      @      4@      @       @      �?      (@              @      �?      @      2@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�ThG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hK	hsKqhth)h,K ��h.��R�(KKq��h{�B@         4                     @z����?�           @�@               %                    �?�l5wA��?�            ps@     �?                           �?�'�=z��?�            �l@                                   �?V�a�� �?Z             b@      �?                          �G@��Q��?)             N@2��                          ��$:@��+7��?             G@ '7��  ������������������������       �                      @�/7��         	                 `f�;@�����?             C@ )7��  ������������������������       �r�q��?             @      @
                        �!�I@     ��?             @@     @                          �<@�����H�?             2@     �?������������������������       ��<ݚ�?             "@        ������������������������       �                     "@       @������������������������       �X�Cc�?
             ,@       @                          �J@X�Cc�?
             ,@     �A@������������������������       �                      @      @������������������������       �r�q��?             @Z                                 �?�̨�`<�?1            @U@       ������������������������       �z�G�z�?             $@�                                �@@���Lͩ�?,            �R@                                 5@�nkK�?             G@       ������������������������       �"pc�
�?             &@�      ������������������������       �                    �A@�                                �E@д>��C�?             =@                                 �B@X�Cc�?	             ,@      ������������������������       �      �?              @c      ������������������������       �      �?             @      ������������������������       �        	             .@                                  :@ �#�Ѵ�?9            �U@                                 �3@��2(&�?             6@       ������������������������       �      �?              @V      ������������������������       �        
             ,@J      !       "                   �H@     ��?+             P@      ������������������������       �        "            �I@A      #       $                   @K@$�q-�?	             *@        ������������������������       �z�G�z�?             @�       ������������������������       �                      @v       &       /                    �?���Q8�?4             T@        '       *                    �?���@M^�?             ?@        (       )                    �?z�G�z�?             $@        ������������������������       �r�q��?             @�       ������������������������       �      �?             @�       +       ,                   �:@�G��l��?             5@        ������������������������       �                     @       -       .                   �>@     ��?
             0@        ������������������������       �r�q��?             @-       ������������������������       ����Q��?             $@]       0       3                   �:@Hm_!'1�?            �H@       1       2                 ��[@؇���X�?             <@       ������������������������       �                     3@�       ������������������������       �X�<ݚ�?             "@�       ������������������������       �                     5@�       5       Z                 `f�%@1`�N�?�            y@       6       Q                    �?l ��H|�?�            �p@      7       D                 �{@X�M|H�?�            `k@        8       ?                  ��@`{��T��??            @Y@      9       :                 `f�@     �?)             P@       ������������������������       �      �?             @;      ;       >                   �;@(;L]n�?%             N@       <       =                   �4@�8��8��?             8@       ������������������������       �                      @7      ������������������������       �      �?
             0@G       ������������������������       �                     B@      @       A                    �?���"͏�?            �B@       ������������������������       ��<ݚ�?
             2@�      B       C                    ;@�d�����?             3@      ������������������������       ��8��8��?             (@8       ������������������������       �և���X�?             @8      E       F                 �?�@�1e�3��?H            �]@       ������������������������       �                    �C@-      G       J                   �:@p`q�q��?3            �S@       H       I                 ��Y @(;L]n�?             >@       ������������������������       ��C��2(�?             &@�       ������������������������       �                     3@�       K       N                 ��) @�q��/��?            �H@      L       M                    C@�FVQ&�?            �@@      ������������������������       �                     :@�      ������������������������       �����X�?             @�      O       P                 @Q!@      �?	             0@       ������������������������       �����X�?             @�      ������������������������       ��<ݚ�?             "@�       R       S                    �?�~8�e�?"            �I@       ������������������������       ��<ݚ�?             2@-      T       Y                   �;@r٣����?            �@@      U       X                 ��,#@�LQ�1	�?             7@      V       W                   �4@j���� �?             1@        ������������������������       ����!pc�?             &@y       ������������������������       ��q�q�?             @}       ������������������������       �r�q��?             @�       ������������������������       �                     $@        [       l                 ��Y7@�c��{-�?L            ``@       \       c                    �?�f���?/            �T@        ]       ^                   �4@�G�z��?             D@        ������������������������       ��r����?             .@        _       `                    �?z�G�z�?             9@        ������������������������       �                     @        a       b                    =@      �?
             4@       ������������������������       ��q�q�?             .@        ������������������������       �                     @        d       k                 ���4@8�$�>�?            �E@       e       f                    �?����X�?            �A@        ������������������������       �      �?              @        g       h                    ;@������?             ;@        ������������������������       ��z�G��?             $@        i       j                 @3�/@������?	             1@        ������������������������       ��q�q�?             @        ������������������������       �"pc�
�?             &@        ������������������������       �      �?              @        m       n                    �?     ��?             H@        ������������������������       �      �?             ,@        o       p                    @�IєX�?             A@        ������������������������       �"pc�
�?             &@        ������������������������       �                     7@        �t�bh�h)h,K ��h.��R�(KKqKK��h\�B       �{@     �p@     �a@      e@     �]@      \@     �\@      >@     �C@      5@      A@      (@       @              :@      (@      �?      @      9@      @      0@       @      @       @      "@              "@      @      @      "@               @      @      �?      S@      "@       @       @      Q@      @      F@       @      "@       @     �A@              8@      @      "@      @      @       @      @      @      .@              @     �T@      @      3@      @      @              ,@      �?     �O@             �I@      �?      (@      �?      @               @      7@     �L@      3@      (@       @       @      @      �?      @      �?      &@      $@              @      &@      @      @      �?      @      @      @     �F@      @      8@              3@      @      @              5@     s@      X@     �l@     �D@      i@      3@     @V@      (@     �N@      @      @      �?      M@       @      6@       @       @              ,@       @      B@              <@      "@      ,@      @      ,@      @      &@      �?      @      @     �[@      @     �C@              R@      @      =@      �?      $@      �?      3@             �E@      @      ?@       @      :@              @       @      (@      @      @       @      @       @      =@      6@      @      ,@      9@       @      .@       @      $@      @       @      @       @      @      @      �?      $@              S@     �K@     �B@      G@      6@      2@       @      *@      4@      @      @              .@      @      $@      @      @              .@      <@      $@      9@      @      @      @      4@      @      @      @      *@       @      @       @      "@      @      @     �C@      "@      @      @      @@       @      "@       @      7@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ5�R/hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsK}hth)h,K ��h.��R�(KK}��h{�B@         X                    �?4�<����?�           @�@                                  @��%n��?&           P}@      (@                        @3�4@�ՙ/�?             5@       @������������������������       �                     @��������������������������������       �և���X�?             ,@      @       ?                 ��D:@     8�?            |@     @       >                    �?س��7'�?�            �t@              	                   �0@$	4�}�?�            t@      ,@������������������������       ��q�q�?             "@      @
                        ��@,�T�6�?�            �s@       @                        ���@     ��?             @@      @                           ?@R���Q�?             4@     �?������������������������       �z�G�z�?
             .@        ������������������������       �                     @      @������������������������       ��q�q�?             (@      �?       5                   @A@�d�g��?�            �q@              ,                   �<@�s��2��?�            �k@                              �?�@�8��8��?l             e@                               �?$@���7�?6             V@                                 �?$�q-�?              J@                               ���@@4և���?             ,@       ������������������������       �r�q��?             @�      ������������������������       �                      @�                                 �?�˹�m��?             C@       ������������������������       �$�q-�?             *@�                              ��@HP�s��?             9@      ������������������������       �        
             5@      ������������������������       �      �?             @      ������������������������       �                     B@�                                �2@      �?6             T@       ������������������������       �                     "@V              #                 pf� @D��\��?0            �Q@       !       "                    ;@R�}e�.�?             :@       ������������������������       �z�G�z�?             $@A      ������������������������       �     ��?
             0@�       $       %                    6@��S�ۿ?             �F@        ������������������������       �z�G�z�?             @v       &       +                    �?P���Q�?             D@       '       *                 ���/@�>����?             ;@       (       )                     @���N8�?             5@       ������������������������       �$�q-�?	             *@�       ������������������������       �                      @�       ������������������������       �r�q��?             @$       ������������������������       �        	             *@       -       .                     @D>�Q�?             J@        ������������������������       ��z�G��?             $@-       /       4                   @@@؇���X�?             E@       0       3                 @3�@�n`���?             ?@       1       2                 �&B@�d�����?             3@        ������������������������       ������H�?             "@�       ������������������������       ����Q��?             $@�       ������������������������       ��8��8��?             (@�       ������������������������       �                     &@�       6       =                   �*@P���Q�?"             N@      7       8                 �?�@�˹�m��?             C@        ������������������������       �                     4@`      9       :                   �B@r�q��?             2@       ������������������������       �                     @;      ;       <                 `f'@      �?	             (@      ������������������������       ����Q��?             @I      ������������������������       �؇���X�?             @7      ������������������������       �        
             6@G       ������������������������       �      �?              @      @       U                     �?��5Վ3�?O            �]@      A       D                   �;@�û��|�?9             W@       B       C                    7@j���� �?	             1@      ������������������������       �      �?              @8       ������������������������       ��<ݚ�?             "@8      E       P                    �?.�W����?0            �R@      F       O                    �?��V#�?            �E@      G       J                    �?p�ݯ��?             C@       H       I                    ?@����X�?	             ,@       ������������������������       �                      @�       ������������������������       ��q�q�?             @�       K       N                   �>@�q�q�?             8@      L       M                   �I@�q�q�?
             .@      ������������������������       �؇���X�?             @�      ������������������������       �      �?              @�      ������������������������       �                     "@�      ������������������������       �                     @�      Q       R                    �?      �?             @@        ������������������������       �      �?              @      S       T                   �D@�q�q�?             8@       ������������������������       �և���X�?             ,@%      ������������������������       �                     $@g      V       W                    �?�����H�?             ;@        ������������������������       �      �?             @y       ������������������������       �                     5@}       Y       f                     @d�� z�?�            `n@       Z       c                  "�b@P�� �?Q            @`@       [       `                   �H@h�����?F             \@       \       _                    6@`Ql�R�?;            �W@        ]       ^                   �;@���}<S�?             7@        ������������������������       ��<ݚ�?             "@        ������������������������       �        	             ,@        ������������������������       �        ,            �Q@        a       b                    �?�����H�?             2@       ������������������������       �      �?              @        ������������������������       �                     $@        d       e                 `D�c@�E��ӭ�?             2@        ������������������������       �      �?              @        ������������������������       �                     $@        g       z                    @+Y���?G            @\@       h       m                    �?     ��?<             X@        i       l                  S�-@��i#[�?             E@       j       k                   �0@�P�*�?             ?@        ������������������������       �r�q��?             @        ������������������������       ��q�����?             9@        ������������������������       �                     &@        n       y                    @�5��?#             K@       o       v                    �?Tt�ó��?            �H@       p       q                   �4@<=�,S��?            �A@        ������������������������       �z�G�z�?             $@        r       s                   #@� �	��?             9@        ������������������������       �      �?             (@        t       u                 ���*@�n_Y�K�?	             *@        ������������������������       ��q�q�?             @        ������������������������       �և���X�?             @        w       x                 `fF5@X�Cc�?	             ,@       ������������������������       �      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     @        {       |                   �0@�t����?             1@       ������������������������       �                     &@        ������������������������       ��q�q�?             @        �t�bh�h)h,K ��h.��R�(KK}KK��h\�B�        |@     �p@     �w@     �V@       @      *@              @       @      @     0w@     @S@     0r@      C@     �q@      B@      @      @     pq@     �@@      9@      @      1@      @      (@      @      @               @      @     �o@      :@     �h@      7@     @c@      ,@      U@      @      H@      @      *@      �?      @      �?       @             �A@      @      (@      �?      7@       @      5@               @       @      B@             �Q@      $@      "@             �N@      $@      3@      @       @       @      &@      @      E@      @      @      �?      C@       @      9@       @      4@      �?      (@      �?       @              @      �?      *@             �E@      "@      @      @      B@      @      9@      @      ,@      @       @      �?      @      @      &@      �?      &@             �L@      @     �A@      @      4@              .@      @      @              "@      @      @       @      @      �?      6@              @       @      T@     �C@      L@      B@      @      $@      @      @       @      @     �H@      :@      =@      ,@      8@      ,@      $@      @       @               @      @      ,@      $@      @      $@      �?      @      @      @      "@              @              4@      (@      @      @      0@       @      @       @      $@              8@      @      @      @      5@             @Q@     �e@      "@     @^@      @      [@       @      W@       @      5@       @      @              ,@             �Q@       @      0@       @      @              $@      @      *@      @      @              $@      N@     �J@     �F@     �I@      *@      =@      *@      2@      �?      @      (@      *@              &@      @@      6@      ;@      6@      6@      *@       @       @      ,@      &@      "@      @      @       @       @      @      @      @      @      "@      �?      @      @       @      @              .@       @      &@              @       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hG?�      hNhJ�%hG        hNhG        hBKhCKhDh)h,K ��h.��R�(KK��h\�C              �?�t�bhPhahKC       ���R�heKhfhiKh)h,K ��h.��R�(KK��hK�C       �t�bK��R�}�(hKhsKwhth)h,K ��h.��R�(KKw��h{�B�         .                     @
Ϛ����?�           @�@               !                    �?�p/����?�            �r@                                   �?u-�KW�?p            �e@     @                        Ј�U@P*L�9�?<             V@     @                          �;@<ݚ�?1             R@      @������������������������       �X�<ݚ�?             "@      @                          �B@Z���c��?,            �O@      @       	                   �G@">�֕�?            �A@     $@������������������������       ��GN�z�?             6@        
                          �L@��
ц��?	             *@      I@������������������������       �r�q��?             @      8@������������������������       �؇���X�?             @      F@                         x#J@@4և���?             <@      C@������������������������       �                     &@      6@                        Ј@S@�t����?             1@      �?������������������������       �      �?              @      @������������������������       �                     "@Z                                �D@      �?             0@      ������������������������       ��<ݚ�?             "@�      ������������������������       �և���X�?             @w                                 ,@�:���?4            �U@                                �7@ �h�7W�?            �J@       ������������������������       �؇���X�?             @�                                �@@�nkK�?             G@       ������������������������       �                     9@�                              `f�)@�����?             5@       ������������������������       �                     "@      ������������������������       �r�q��?             (@                                 "@H�V�e��?             A@       ������������������������       �                     @(                                 �@@h�����?             <@       ������������������������       �ףp=
�?             $@J      ������������������������       �        
             2@3      "       +                  "�b@`Jj��?W             _@      #       &                   �;@ 7���B�?M             [@        $       %                   �7@��S�ۿ?            �F@       ������������������������       �                     ?@v       ������������������������       �d}h���?             ,@j       '       *                     �? ������?0            �O@       (       )                   �H@      �?             @@       ������������������������       �                     6@�       ������������������������       �ףp=
�?             $@�       ������������������������       �                     ?@$       ,       -                    �?      �?
             0@       ������������������������       �                     $@       ������������������������       ��q�q�?             @-       /       `                 `�X.@2�����?           �y@       0       ]                    �?���_�?�             s@       1       R                    �?�)Kj	�?�            �q@       2       O                   @@@=�J�C�?�            �m@       3       N                    �?,sI�v�?o            �f@       4       9                    �?��㨇,�?j            �e@        5       6                 ���@@4և���?             E@        ������������������������       �                     $@      7       8                   �:@     ��?             @@        ������������������������       ��q�q�?             @`      ������������������������       � ��WV�?             :@:      :       A                   �7@ ����?O            ``@       ;       <                 �?�@l�b�G��?             �L@       ������������������������       �                     >@I      =       @                   �3@PN��T'�?             ;@      >       ?                 ��Y @������?
             .@        ������������������������       ��q�q�?             @      ������������������������       �                     "@!      ������������������������       �                     (@�      B       E                 ��]@��A��?/            �R@       C       D                 pf�@ҳ�wY;�?             1@       ������������������������       �z�G�z�?             $@8      ������������������������       �և���X�?             @      F       K                 ��) @���5��?$            �L@      G       H                 �?�@�7��?            �C@      ������������������������       �                     3@�      I       J                   �<@ףp=
�?
             4@       ������������������������       �                     (@�       ������������������������       �      �?              @v      L       M                 0S%"@�E��ӭ�?             2@       ������������������������       ��q�q�?             "@�      ������������������������       ��<ݚ�?             "@�      ������������������������       �����X�?             @�      P       Q                 �?�@P����?#            �M@      ������������������������       �                     A@�       ������������������������       �`2U0*��?             9@      S       \                 pF @��C���?            �G@      T       Y                   �9@J�8���?             =@      U       X                   �5@��S���?             .@      V       W                  s�@�q�q�?             "@        ������������������������       �                     @y       ������������������������       �      �?             @}       ������������������������       �r�q��?             @�       Z       [                 �Y5@؇���X�?	             ,@       ������������������������       �����X�?             @        ������������������������       �                     @        ������������������������       �        
             2@        ^       _                    �?���Q��?             4@        ������������������������       ����!pc�?             &@        ������������������������       �X�<ݚ�?             "@        a       r                    @r�0?��?E            �Z@       b       c                    �?�):u��?1            @S@        ������������������������       �                     *@        d       m                    �?     x�?)             P@       e       l                   @@@�d�����?             C@       f       g                    �?�q�q�?             >@        ������������������������       �      �?              @        h       k                 �T)D@8�A�0��?             6@       i       j                   �2@z�G�z�?
             .@        ������������������������       �      �?             @        ������������������������       �                     "@        ������������������������       �؇���X�?             @        ������������������������       �                      @        n       q                   �<@      �?             :@       o       p                    :@�q�q�?	             .@        ������������������������       �և���X�?             @        ������������������������       �      �?              @        ������������������������       ����!pc�?             &@        s       t                    �?ףp=
�?             >@        ������������������������       �                     ,@        u       v                 pf�C@     ��?             0@        ������������������������       �և���X�?             @        ������������������������       �                     "@        �t�bh�h)h,K ��h.��R�(KKwKK��h\�Bp       `}@     @n@     @b@      c@     @a@     �B@     �N@      ;@     �K@      1@      @      @      I@      *@      8@      &@      1@      @      @      @      �?      @      @      �?      :@       @      &@              .@       @      @       @      "@              @      $@       @      @      @      @     @S@      $@      I@      @      @      �?      F@       @      9@              3@       @      "@              $@       @      ;@      @              @      ;@      �?      "@      �?      2@               @      ]@      @      Z@      @      E@              ?@      @      &@      �?      O@      �?      ?@              6@      �?      "@              ?@      @      (@              $@      @       @     @t@     @V@      p@      I@     �n@      E@      k@      7@     �c@      6@      c@      4@     �C@      @      $@              =@      @      @       @      9@      �?     �\@      1@     �J@      @      >@              7@      @      &@      @       @      @      "@              (@             �N@      *@      &@      @       @       @      @      @      I@      @     �B@       @      3@              2@       @      (@              @       @      *@      @      @      @      @       @      @       @      M@      �?      A@              8@      �?      <@      3@      $@      3@       @      @      @      @              @      @      �?      @      �?       @      (@       @      @              @      2@              (@       @       @      @      @      @      Q@     �C@     �D@      B@              *@     �D@      7@      <@      $@      4@      $@      @      �?      *@      "@      (@      @      @      @      "@              �?      @       @              *@      *@      @      $@      @      @      �?      @       @      @      ;@      @      ,@              *@      @      @      @      "@        �t�bubhhubehhub.